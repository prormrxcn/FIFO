magic
tech sky130A
magscale 1 2
timestamp 1755446084
<< checkpaint >>
rect -1260 8876 34234 36378
rect -2590 372 34234 8876
rect -1260 -1260 34234 372
<< viali >>
rect 19441 32521 19475 32555
rect 24961 32521 24995 32555
rect 1409 32385 1443 32419
rect 7205 32385 7239 32419
rect 13001 32385 13035 32419
rect 19349 32385 19383 32419
rect 24685 32385 24719 32419
rect 30389 32385 30423 32419
rect 1593 32249 1627 32283
rect 7389 32181 7423 32215
rect 13185 32181 13219 32215
rect 30573 32181 30607 32215
rect 19901 31773 19935 31807
rect 19257 31637 19291 31671
rect 13553 31433 13587 31467
rect 15577 31433 15611 31467
rect 17693 31365 17727 31399
rect 18705 31365 18739 31399
rect 11989 31297 12023 31331
rect 12357 31297 12391 31331
rect 13277 31297 13311 31331
rect 13737 31297 13771 31331
rect 16957 31297 16991 31331
rect 17049 31297 17083 31331
rect 17141 31297 17175 31331
rect 17325 31297 17359 31331
rect 17417 31297 17451 31331
rect 17509 31297 17543 31331
rect 17785 31297 17819 31331
rect 17877 31297 17911 31331
rect 18061 31297 18095 31331
rect 12081 31229 12115 31263
rect 12909 31229 12943 31263
rect 13829 31229 13863 31263
rect 14105 31229 14139 31263
rect 18429 31229 18463 31263
rect 17693 31161 17727 31195
rect 18061 31161 18095 31195
rect 20177 31161 20211 31195
rect 11621 31093 11655 31127
rect 13185 31093 13219 31127
rect 16865 31093 16899 31127
rect 17325 31093 17359 31127
rect 13737 30889 13771 30923
rect 14841 30889 14875 30923
rect 18429 30889 18463 30923
rect 21017 30889 21051 30923
rect 12541 30821 12575 30855
rect 18337 30821 18371 30855
rect 11069 30753 11103 30787
rect 15485 30753 15519 30787
rect 21281 30753 21315 30787
rect 1409 30685 1443 30719
rect 10793 30685 10827 30719
rect 13185 30685 13219 30719
rect 13553 30685 13587 30719
rect 14289 30685 14323 30719
rect 14749 30685 14783 30719
rect 17969 30685 18003 30719
rect 18153 30685 18187 30719
rect 18337 30685 18371 30719
rect 19073 30685 19107 30719
rect 19257 30685 19291 30719
rect 13369 30617 13403 30651
rect 13461 30617 13495 30651
rect 15761 30617 15795 30651
rect 1593 30549 1627 30583
rect 14197 30549 14231 30583
rect 17233 30549 17267 30583
rect 17417 30549 17451 30583
rect 15669 30345 15703 30379
rect 15853 30345 15887 30379
rect 14749 30277 14783 30311
rect 19073 30277 19107 30311
rect 11897 30209 11931 30243
rect 12633 30209 12667 30243
rect 13921 30209 13955 30243
rect 14933 30209 14967 30243
rect 15794 30209 15828 30243
rect 16221 30209 16255 30243
rect 17601 30209 17635 30243
rect 17877 30209 17911 30243
rect 18521 30209 18555 30243
rect 15117 30141 15151 30175
rect 16313 30141 16347 30175
rect 16773 30141 16807 30175
rect 17969 30141 18003 30175
rect 18245 30141 18279 30175
rect 18797 30141 18831 30175
rect 13553 30005 13587 30039
rect 14013 30005 14047 30039
rect 18613 30005 18647 30039
rect 20545 30005 20579 30039
rect 13921 29801 13955 29835
rect 14105 29801 14139 29835
rect 16221 29801 16255 29835
rect 16681 29801 16715 29835
rect 16865 29801 16899 29835
rect 19441 29801 19475 29835
rect 19717 29801 19751 29835
rect 15669 29733 15703 29767
rect 13001 29665 13035 29699
rect 17509 29665 17543 29699
rect 13369 29597 13403 29631
rect 13461 29597 13495 29631
rect 13553 29597 13587 29631
rect 13737 29597 13771 29631
rect 14289 29597 14323 29631
rect 14473 29597 14507 29631
rect 15485 29597 15519 29631
rect 16405 29597 16439 29631
rect 16589 29597 16623 29631
rect 17693 29597 17727 29631
rect 17877 29597 17911 29631
rect 19349 29597 19383 29631
rect 19625 29597 19659 29631
rect 17049 29529 17083 29563
rect 13277 29461 13311 29495
rect 16839 29461 16873 29495
rect 14565 29121 14599 29155
rect 14749 28985 14783 29019
rect 12357 28713 12391 28747
rect 8493 28509 8527 28543
rect 8953 28509 8987 28543
rect 10609 28509 10643 28543
rect 14381 28509 14415 28543
rect 9198 28441 9232 28475
rect 10885 28441 10919 28475
rect 14289 28441 14323 28475
rect 14657 28441 14691 28475
rect 8677 28373 8711 28407
rect 10333 28373 10367 28407
rect 14105 28373 14139 28407
rect 14473 28373 14507 28407
rect 8769 28169 8803 28203
rect 13737 28169 13771 28203
rect 13829 28169 13863 28203
rect 14933 28169 14967 28203
rect 14841 28101 14875 28135
rect 16957 28101 16991 28135
rect 9137 28033 9171 28067
rect 9781 28033 9815 28067
rect 10885 28033 10919 28067
rect 11621 28033 11655 28067
rect 12173 28033 12207 28067
rect 13369 28033 13403 28067
rect 13645 28033 13679 28067
rect 14289 28033 14323 28067
rect 14381 28033 14415 28067
rect 14473 28033 14507 28067
rect 16681 28033 16715 28067
rect 16865 28033 16899 28067
rect 17877 28033 17911 28067
rect 20361 28033 20395 28067
rect 23397 28033 23431 28067
rect 26617 28033 26651 28067
rect 9229 27965 9263 27999
rect 9321 27965 9355 27999
rect 10333 27965 10367 27999
rect 10517 27965 10551 27999
rect 10793 27965 10827 27999
rect 13185 27965 13219 27999
rect 16497 27965 16531 27999
rect 18061 27965 18095 27999
rect 20269 27965 20303 27999
rect 14013 27897 14047 27931
rect 14657 27897 14691 27931
rect 16221 27897 16255 27931
rect 17325 27897 17359 27931
rect 20729 27897 20763 27931
rect 13461 27829 13495 27863
rect 14105 27829 14139 27863
rect 16037 27829 16071 27863
rect 16681 27829 16715 27863
rect 17417 27829 17451 27863
rect 17693 27829 17727 27863
rect 23213 27829 23247 27863
rect 26433 27829 26467 27863
rect 16773 27557 16807 27591
rect 17417 27557 17451 27591
rect 19809 27557 19843 27591
rect 20729 27557 20763 27591
rect 14724 27489 14758 27523
rect 19349 27489 19383 27523
rect 19993 27489 20027 27523
rect 9045 27421 9079 27455
rect 11069 27421 11103 27455
rect 13829 27421 13863 27455
rect 14933 27421 14967 27455
rect 15209 27421 15243 27455
rect 16129 27421 16163 27455
rect 16614 27421 16648 27455
rect 17785 27421 17819 27455
rect 18061 27421 18095 27455
rect 18705 27421 18739 27455
rect 18981 27421 19015 27455
rect 19441 27421 19475 27455
rect 20085 27421 20119 27455
rect 21005 27421 21039 27455
rect 22845 27421 22879 27455
rect 23112 27421 23146 27455
rect 24961 27421 24995 27455
rect 26065 27421 26099 27455
rect 26332 27421 26366 27455
rect 28089 27421 28123 27455
rect 7113 27353 7147 27387
rect 7481 27353 7515 27387
rect 9312 27353 9346 27387
rect 13461 27353 13495 27387
rect 17693 27353 17727 27387
rect 18337 27353 18371 27387
rect 21281 27353 21315 27387
rect 10425 27285 10459 27319
rect 10517 27285 10551 27319
rect 14565 27285 14599 27319
rect 14841 27285 14875 27319
rect 16405 27285 16439 27319
rect 16497 27285 16531 27319
rect 17601 27285 17635 27319
rect 17969 27285 18003 27319
rect 18705 27285 18739 27319
rect 20453 27285 20487 27319
rect 20913 27285 20947 27319
rect 21097 27285 21131 27319
rect 24225 27285 24259 27319
rect 24409 27285 24443 27319
rect 27445 27285 27479 27319
rect 27537 27285 27571 27319
rect 9229 27081 9263 27115
rect 9873 27081 9907 27115
rect 15025 27081 15059 27115
rect 17049 27081 17083 27115
rect 17233 27081 17267 27115
rect 18337 27081 18371 27115
rect 18429 27081 18463 27115
rect 20913 27081 20947 27115
rect 23305 27081 23339 27115
rect 23673 27081 23707 27115
rect 26985 27081 27019 27115
rect 27353 27081 27387 27115
rect 28549 27081 28583 27115
rect 8125 27013 8159 27047
rect 15234 27013 15268 27047
rect 16338 27013 16372 27047
rect 16681 27013 16715 27047
rect 17601 27013 17635 27047
rect 19441 27013 19475 27047
rect 25688 27013 25722 27047
rect 7757 26945 7791 26979
rect 9413 26945 9447 26979
rect 13369 26945 13403 26979
rect 13737 26945 13771 26979
rect 14381 26945 14415 26979
rect 16129 26945 16163 26979
rect 16865 26945 16899 26979
rect 16957 26945 16991 26979
rect 17693 26945 17727 26979
rect 17810 26945 17844 26979
rect 18797 26945 18831 26979
rect 20545 26945 20579 26979
rect 23765 26945 23799 26979
rect 27445 26945 27479 26979
rect 28733 26945 28767 26979
rect 7389 26877 7423 26911
rect 9965 26877 9999 26911
rect 10149 26877 10183 26911
rect 12541 26877 12575 26911
rect 13921 26877 13955 26911
rect 14289 26877 14323 26911
rect 14776 26877 14810 26911
rect 15117 26877 15151 26911
rect 15853 26877 15887 26911
rect 16221 26877 16255 26911
rect 17325 26877 17359 26911
rect 18061 26877 18095 26911
rect 18546 26877 18580 26911
rect 19073 26877 19107 26911
rect 20453 26877 20487 26911
rect 23949 26877 23983 26911
rect 25421 26877 25455 26911
rect 27537 26877 27571 26911
rect 28365 26877 28399 26911
rect 9505 26809 9539 26843
rect 12817 26809 12851 26843
rect 16497 26809 16531 26843
rect 17969 26809 18003 26843
rect 26801 26809 26835 26843
rect 6745 26741 6779 26775
rect 14565 26741 14599 26775
rect 15393 26741 15427 26775
rect 18705 26741 18739 26775
rect 19717 26741 19751 26775
rect 27813 26741 27847 26775
rect 6653 26537 6687 26571
rect 15301 26537 15335 26571
rect 18153 26537 18187 26571
rect 27997 26537 28031 26571
rect 8125 26469 8159 26503
rect 15853 26469 15887 26503
rect 17509 26469 17543 26503
rect 9505 26401 9539 26435
rect 14841 26401 14875 26435
rect 16865 26401 16899 26435
rect 17141 26401 17175 26435
rect 17233 26401 17267 26435
rect 25789 26401 25823 26435
rect 27445 26401 27479 26435
rect 5273 26333 5307 26367
rect 6745 26333 6779 26367
rect 13369 26333 13403 26367
rect 13921 26333 13955 26367
rect 14565 26333 14599 26367
rect 14933 26333 14967 26367
rect 17877 26333 17911 26367
rect 18245 26333 18279 26367
rect 19349 26333 19383 26367
rect 19717 26333 19751 26367
rect 23489 26333 23523 26367
rect 23673 26333 23707 26367
rect 24961 26333 24995 26367
rect 27629 26333 27663 26367
rect 5540 26265 5574 26299
rect 7012 26265 7046 26299
rect 13093 26265 13127 26299
rect 13645 26265 13679 26299
rect 15050 26265 15084 26299
rect 15485 26265 15519 26299
rect 15577 26265 15611 26299
rect 15669 26265 15703 26299
rect 17350 26265 17384 26299
rect 17601 26265 17635 26299
rect 17969 26265 18003 26299
rect 18521 26265 18555 26299
rect 19901 26265 19935 26299
rect 26056 26265 26090 26299
rect 31125 26265 31159 26299
rect 31493 26265 31527 26299
rect 8953 26197 8987 26231
rect 15209 26197 15243 26231
rect 17785 26197 17819 26231
rect 20177 26197 20211 26231
rect 23305 26197 23339 26231
rect 23857 26197 23891 26231
rect 24409 26197 24443 26231
rect 27169 26197 27203 26231
rect 27537 26197 27571 26231
rect 6745 25993 6779 26027
rect 7297 25993 7331 26027
rect 7573 25993 7607 26027
rect 7849 25993 7883 26027
rect 8217 25993 8251 26027
rect 14105 25993 14139 26027
rect 14289 25993 14323 26027
rect 4905 25925 4939 25959
rect 6653 25925 6687 25959
rect 9965 25925 9999 25959
rect 14381 25925 14415 25959
rect 15117 25925 15151 25959
rect 15393 25925 15427 25959
rect 19533 25925 19567 25959
rect 29193 25925 29227 25959
rect 4537 25857 4571 25891
rect 4997 25857 5031 25891
rect 5457 25857 5491 25891
rect 7481 25857 7515 25891
rect 7757 25857 7791 25891
rect 9689 25857 9723 25891
rect 9837 25857 9871 25891
rect 10057 25857 10091 25891
rect 10154 25857 10188 25891
rect 14473 25857 14507 25891
rect 18889 25857 18923 25891
rect 23204 25857 23238 25891
rect 24409 25857 24443 25891
rect 24665 25857 24699 25891
rect 26433 25857 26467 25891
rect 26985 25857 27019 25891
rect 4813 25789 4847 25823
rect 6009 25789 6043 25823
rect 6561 25789 6595 25823
rect 8309 25789 8343 25823
rect 8493 25789 8527 25823
rect 19165 25789 19199 25823
rect 22937 25789 22971 25823
rect 26525 25789 26559 25823
rect 26709 25789 26743 25823
rect 27629 25789 27663 25823
rect 7113 25721 7147 25755
rect 14657 25721 14691 25755
rect 24317 25721 24351 25755
rect 29377 25721 29411 25755
rect 4353 25653 4387 25687
rect 5365 25653 5399 25687
rect 10333 25653 10367 25687
rect 14841 25653 14875 25687
rect 15669 25653 15703 25687
rect 19809 25653 19843 25687
rect 25789 25653 25823 25687
rect 26065 25653 26099 25687
rect 5457 25449 5491 25483
rect 9689 25449 9723 25483
rect 23489 25449 23523 25483
rect 24409 25449 24443 25483
rect 5365 25381 5399 25415
rect 12173 25381 12207 25415
rect 3985 25313 4019 25347
rect 5917 25313 5951 25347
rect 6009 25313 6043 25347
rect 12817 25313 12851 25347
rect 24041 25313 24075 25347
rect 25053 25313 25087 25347
rect 25881 25313 25915 25347
rect 6929 25245 6963 25279
rect 7297 25245 7331 25279
rect 9505 25245 9539 25279
rect 9873 25245 9907 25279
rect 9965 25245 9999 25279
rect 10241 25245 10275 25279
rect 10793 25245 10827 25279
rect 19441 25245 19475 25279
rect 20453 25245 20487 25279
rect 23857 25245 23891 25279
rect 26249 25245 26283 25279
rect 4252 25177 4286 25211
rect 5825 25177 5859 25211
rect 6285 25177 6319 25211
rect 7564 25177 7598 25211
rect 10057 25177 10091 25211
rect 11060 25177 11094 25211
rect 23949 25177 23983 25211
rect 24777 25177 24811 25211
rect 25329 25177 25363 25211
rect 8677 25109 8711 25143
rect 8953 25109 8987 25143
rect 12265 25109 12299 25143
rect 19349 25109 19383 25143
rect 20637 25109 20671 25143
rect 24869 25109 24903 25143
rect 26065 25109 26099 25143
rect 5365 24905 5399 24939
rect 7757 24905 7791 24939
rect 8401 24905 8435 24939
rect 11161 24905 11195 24939
rect 11897 24905 11931 24939
rect 19901 24905 19935 24939
rect 29653 24905 29687 24939
rect 4160 24837 4194 24871
rect 24501 24837 24535 24871
rect 29561 24837 29595 24871
rect 30297 24837 30331 24871
rect 3893 24769 3927 24803
rect 5549 24769 5583 24803
rect 7941 24769 7975 24803
rect 10885 24769 10919 24803
rect 10977 24769 11011 24803
rect 11345 24769 11379 24803
rect 11989 24769 12023 24803
rect 14013 24769 14047 24803
rect 20085 24769 20119 24803
rect 24225 24769 24259 24803
rect 24409 24769 24443 24803
rect 24593 24769 24627 24803
rect 25421 24769 25455 24803
rect 25605 24769 25639 24803
rect 25697 24769 25731 24803
rect 25789 24769 25823 24803
rect 27169 24769 27203 24803
rect 27261 24769 27295 24803
rect 27353 24769 27387 24803
rect 27537 24769 27571 24803
rect 30021 24769 30055 24803
rect 1409 24701 1443 24735
rect 1685 24701 1719 24735
rect 8493 24701 8527 24735
rect 8585 24701 8619 24735
rect 8953 24701 8987 24735
rect 9229 24701 9263 24735
rect 12173 24701 12207 24735
rect 13737 24701 13771 24735
rect 18153 24701 18187 24735
rect 18429 24701 18463 24735
rect 28549 24701 28583 24735
rect 29745 24701 29779 24735
rect 30849 24701 30883 24735
rect 5273 24633 5307 24667
rect 8033 24633 8067 24667
rect 10701 24633 10735 24667
rect 11529 24633 11563 24667
rect 13921 24633 13955 24667
rect 13829 24565 13863 24599
rect 20177 24565 20211 24599
rect 24777 24565 24811 24599
rect 25973 24565 26007 24599
rect 26985 24565 27019 24599
rect 29101 24565 29135 24599
rect 29193 24565 29227 24599
rect 30205 24565 30239 24599
rect 9321 24361 9355 24395
rect 16681 24361 16715 24395
rect 18889 24361 18923 24395
rect 20085 24361 20119 24395
rect 25973 24361 26007 24395
rect 29377 24361 29411 24395
rect 6101 24293 6135 24327
rect 8493 24293 8527 24327
rect 11437 24293 11471 24327
rect 26249 24293 26283 24327
rect 10333 24225 10367 24259
rect 11805 24225 11839 24259
rect 16313 24225 16347 24259
rect 19926 24225 19960 24259
rect 20545 24225 20579 24259
rect 21373 24225 21407 24259
rect 25973 24225 26007 24259
rect 28825 24225 28859 24259
rect 28917 24225 28951 24259
rect 5549 24157 5583 24191
rect 5917 24157 5951 24191
rect 8033 24157 8067 24191
rect 8309 24157 8343 24191
rect 9505 24157 9539 24191
rect 10057 24157 10091 24191
rect 11253 24157 11287 24191
rect 11345 24157 11379 24191
rect 11529 24157 11563 24191
rect 13461 24157 13495 24191
rect 14657 24157 14691 24191
rect 15025 24157 15059 24191
rect 16405 24157 16439 24191
rect 18981 24157 19015 24191
rect 19441 24157 19475 24191
rect 20269 24157 20303 24191
rect 20361 24157 20395 24191
rect 20453 24157 20487 24191
rect 21465 24157 21499 24191
rect 21557 24157 21591 24191
rect 21649 24157 21683 24191
rect 22937 24157 22971 24191
rect 23213 24157 23247 24191
rect 25789 24157 25823 24191
rect 26065 24157 26099 24191
rect 28365 24157 28399 24191
rect 29561 24157 29595 24191
rect 5733 24089 5767 24123
rect 5825 24089 5859 24123
rect 8125 24089 8159 24123
rect 11989 24089 12023 24123
rect 12173 24089 12207 24123
rect 13277 24089 13311 24123
rect 13829 24089 13863 24123
rect 14197 24089 14231 24123
rect 20729 24089 20763 24123
rect 21833 24089 21867 24123
rect 24961 24089 24995 24123
rect 25145 24089 25179 24123
rect 29009 24089 29043 24123
rect 29806 24089 29840 24123
rect 9689 24021 9723 24055
rect 10149 24021 10183 24055
rect 11713 24021 11747 24055
rect 13553 24021 13587 24055
rect 13645 24021 13679 24055
rect 14289 24021 14323 24055
rect 14841 24021 14875 24055
rect 15117 24021 15151 24055
rect 19717 24021 19751 24055
rect 19809 24021 19843 24055
rect 28549 24021 28583 24055
rect 30941 24021 30975 24055
rect 15945 23817 15979 23851
rect 19257 23817 19291 23851
rect 28457 23817 28491 23851
rect 13645 23749 13679 23783
rect 13737 23749 13771 23783
rect 14565 23749 14599 23783
rect 15577 23749 15611 23783
rect 19625 23749 19659 23783
rect 20269 23749 20303 23783
rect 20637 23749 20671 23783
rect 24777 23749 24811 23783
rect 13185 23681 13219 23715
rect 13277 23681 13311 23715
rect 14473 23681 14507 23715
rect 15117 23681 15151 23715
rect 15301 23681 15335 23715
rect 15761 23681 15795 23715
rect 19441 23681 19475 23715
rect 20085 23681 20119 23715
rect 20177 23681 20211 23715
rect 21097 23681 21131 23715
rect 21189 23681 21223 23715
rect 23213 23681 23247 23715
rect 26433 23681 26467 23715
rect 28365 23681 28399 23715
rect 28636 23681 28670 23715
rect 28733 23681 28767 23715
rect 28825 23681 28859 23715
rect 29008 23681 29042 23715
rect 29101 23681 29135 23715
rect 30306 23681 30340 23715
rect 30573 23681 30607 23715
rect 12725 23613 12759 23647
rect 14013 23613 14047 23647
rect 14105 23613 14139 23647
rect 15025 23613 15059 23647
rect 19717 23613 19751 23647
rect 20729 23613 20763 23647
rect 21649 23613 21683 23647
rect 23489 23613 23523 23647
rect 27997 23613 28031 23647
rect 24961 23545 24995 23579
rect 29193 23545 29227 23579
rect 15209 23477 15243 23511
rect 15485 23477 15519 23511
rect 26249 23477 26283 23511
rect 27445 23477 27479 23511
rect 28181 23477 28215 23511
rect 27353 23273 27387 23307
rect 14243 23205 14277 23239
rect 14381 23205 14415 23239
rect 15117 23205 15151 23239
rect 13001 23137 13035 23171
rect 14473 23137 14507 23171
rect 19441 23137 19475 23171
rect 25973 23137 26007 23171
rect 4169 23069 4203 23103
rect 5825 23069 5859 23103
rect 6009 23069 6043 23103
rect 6377 23069 6411 23103
rect 9505 23069 9539 23103
rect 12909 23069 12943 23103
rect 13369 23069 13403 23103
rect 13461 23069 13495 23103
rect 14933 23069 14967 23103
rect 15117 23069 15151 23103
rect 15301 23069 15335 23103
rect 15485 23069 15519 23103
rect 15669 23069 15703 23103
rect 16313 23069 16347 23103
rect 18337 23069 18371 23103
rect 18613 23069 18647 23103
rect 18797 23069 18831 23103
rect 19901 23069 19935 23103
rect 19993 23069 20027 23103
rect 20453 23069 20487 23103
rect 20637 23069 20671 23103
rect 21097 23069 21131 23103
rect 21189 23069 21223 23103
rect 21833 23069 21867 23103
rect 22385 23069 22419 23103
rect 22845 23069 22879 23103
rect 23673 23069 23707 23103
rect 24777 23069 24811 23103
rect 27537 23069 27571 23103
rect 6193 23001 6227 23035
rect 6285 23001 6319 23035
rect 13553 23001 13587 23035
rect 14105 23001 14139 23035
rect 15577 23001 15611 23035
rect 16589 23001 16623 23035
rect 20361 23001 20395 23035
rect 21557 23001 21591 23035
rect 21649 23001 21683 23035
rect 22293 23001 22327 23035
rect 22753 23001 22787 23035
rect 26240 23001 26274 23035
rect 27804 23001 27838 23035
rect 3985 22933 4019 22967
rect 5273 22933 5307 22967
rect 6561 22933 6595 22967
rect 8953 22933 8987 22967
rect 14749 22933 14783 22967
rect 15853 22933 15887 22967
rect 18521 22933 18555 22967
rect 18981 22933 19015 22967
rect 23489 22933 23523 22967
rect 25421 22933 25455 22967
rect 28917 22933 28951 22967
rect 3525 22729 3559 22763
rect 4997 22729 5031 22763
rect 5457 22729 5491 22763
rect 7941 22729 7975 22763
rect 8401 22729 8435 22763
rect 14565 22729 14599 22763
rect 24593 22729 24627 22763
rect 24961 22729 24995 22763
rect 28457 22729 28491 22763
rect 28917 22729 28951 22763
rect 3862 22661 3896 22695
rect 13001 22661 13035 22695
rect 18889 22661 18923 22695
rect 19533 22661 19567 22695
rect 20729 22661 20763 22695
rect 23388 22661 23422 22695
rect 25053 22661 25087 22695
rect 26433 22661 26467 22695
rect 26525 22661 26559 22695
rect 3341 22593 3375 22627
rect 6561 22593 6595 22627
rect 6828 22593 6862 22627
rect 8493 22593 8527 22627
rect 12909 22593 12943 22627
rect 13369 22593 13403 22627
rect 13461 22593 13495 22627
rect 13553 22593 13587 22627
rect 14197 22593 14231 22627
rect 14381 22593 14415 22627
rect 14657 22593 14691 22627
rect 15577 22593 15611 22627
rect 15761 22593 15795 22627
rect 16129 22593 16163 22627
rect 16681 22593 16715 22627
rect 18981 22593 19015 22627
rect 19257 22593 19291 22627
rect 19809 22593 19843 22627
rect 20269 22593 20303 22627
rect 21557 22593 21591 22627
rect 22477 22593 22511 22627
rect 22569 22593 22603 22627
rect 22661 22593 22695 22627
rect 23121 22593 23155 22627
rect 26269 22593 26303 22627
rect 26617 22593 26651 22627
rect 27813 22593 27847 22627
rect 28825 22593 28859 22627
rect 29285 22593 29319 22627
rect 29837 22593 29871 22627
rect 3617 22525 3651 22559
rect 5549 22525 5583 22559
rect 5641 22525 5675 22559
rect 8677 22525 8711 22559
rect 15853 22525 15887 22559
rect 15945 22525 15979 22559
rect 16313 22525 16347 22559
rect 16957 22525 16991 22559
rect 18705 22525 18739 22559
rect 22385 22525 22419 22559
rect 25237 22525 25271 22559
rect 27537 22525 27571 22559
rect 29009 22525 29043 22559
rect 5089 22457 5123 22491
rect 19993 22457 20027 22491
rect 22845 22457 22879 22491
rect 8033 22389 8067 22423
rect 14289 22389 14323 22423
rect 15761 22389 15795 22423
rect 20453 22389 20487 22423
rect 24501 22389 24535 22423
rect 26801 22389 26835 22423
rect 5273 22185 5307 22219
rect 7297 22185 7331 22219
rect 10333 22185 10367 22219
rect 21465 22185 21499 22219
rect 21557 22185 21591 22219
rect 9965 22117 9999 22151
rect 5917 22049 5951 22083
rect 10701 22049 10735 22083
rect 12633 22049 12667 22083
rect 16957 22049 16991 22083
rect 21649 22049 21683 22083
rect 22845 22049 22879 22083
rect 24869 22049 24903 22083
rect 24961 22049 24995 22083
rect 27537 22049 27571 22083
rect 3801 21981 3835 22015
rect 7205 21981 7239 22015
rect 7481 21981 7515 22015
rect 7757 21981 7791 22015
rect 7941 21981 7975 22015
rect 8033 21981 8067 22015
rect 8217 21981 8251 22015
rect 9873 21981 9907 22015
rect 10057 21981 10091 22015
rect 10149 21981 10183 22015
rect 10609 21981 10643 22015
rect 11069 21981 11103 22015
rect 16129 21981 16163 22015
rect 16313 21981 16347 22015
rect 18981 21981 19015 22015
rect 21281 21981 21315 22015
rect 27353 21981 27387 22015
rect 30113 21981 30147 22015
rect 4068 21913 4102 21947
rect 7573 21913 7607 21947
rect 10885 21913 10919 21947
rect 11805 21913 11839 21947
rect 16221 21913 16255 21947
rect 17233 21913 17267 21947
rect 19993 21913 20027 21947
rect 20729 21913 20763 21947
rect 23112 21913 23146 21947
rect 25697 21913 25731 21947
rect 26433 21913 26467 21947
rect 5181 21845 5215 21879
rect 5641 21845 5675 21879
rect 5733 21845 5767 21879
rect 6561 21845 6595 21879
rect 8401 21845 8435 21879
rect 10425 21845 10459 21879
rect 21373 21845 21407 21879
rect 24225 21845 24259 21879
rect 24409 21845 24443 21879
rect 24777 21845 24811 21879
rect 26985 21845 27019 21879
rect 27445 21845 27479 21879
rect 29561 21845 29595 21879
rect 6745 21641 6779 21675
rect 6837 21641 6871 21675
rect 9597 21641 9631 21675
rect 11345 21641 11379 21675
rect 12725 21641 12759 21675
rect 13185 21641 13219 21675
rect 17509 21641 17543 21675
rect 23489 21641 23523 21675
rect 24501 21641 24535 21675
rect 25237 21641 25271 21675
rect 29561 21641 29595 21675
rect 8677 21573 8711 21607
rect 9321 21573 9355 21607
rect 10232 21573 10266 21607
rect 24133 21573 24167 21607
rect 24225 21573 24259 21607
rect 25329 21573 25363 21607
rect 26065 21573 26099 21607
rect 29469 21573 29503 21607
rect 4813 21505 4847 21539
rect 5080 21505 5114 21539
rect 7941 21505 7975 21539
rect 8953 21505 8987 21539
rect 9046 21505 9080 21539
rect 9229 21505 9263 21539
rect 9459 21505 9493 21539
rect 9965 21505 9999 21539
rect 12081 21505 12115 21539
rect 12817 21505 12851 21539
rect 13461 21505 13495 21539
rect 17601 21505 17635 21539
rect 23673 21505 23707 21539
rect 23949 21505 23983 21539
rect 24317 21505 24351 21539
rect 24593 21505 24627 21539
rect 26985 21505 27019 21539
rect 27261 21505 27295 21539
rect 30941 21505 30975 21539
rect 7021 21437 7055 21471
rect 12541 21437 12575 21471
rect 27077 21437 27111 21471
rect 29377 21437 29411 21471
rect 30573 21437 30607 21471
rect 6193 21369 6227 21403
rect 29929 21369 29963 21403
rect 6377 21301 6411 21335
rect 11529 21301 11563 21335
rect 13277 21301 13311 21335
rect 26985 21301 27019 21335
rect 27445 21301 27479 21335
rect 30021 21301 30055 21335
rect 30757 21301 30791 21335
rect 5457 21097 5491 21131
rect 6193 21097 6227 21131
rect 8953 21097 8987 21131
rect 10609 21097 10643 21131
rect 26617 21097 26651 21131
rect 28273 21097 28307 21131
rect 29561 21097 29595 21131
rect 29377 21029 29411 21063
rect 6101 20961 6135 20995
rect 9597 20961 9631 20995
rect 11161 20961 11195 20995
rect 27537 20961 27571 20995
rect 28825 20961 28859 20995
rect 6377 20893 6411 20927
rect 8502 20893 8536 20927
rect 8769 20893 8803 20927
rect 10977 20893 11011 20927
rect 12173 20893 12207 20927
rect 14289 20893 14323 20927
rect 25881 20893 25915 20927
rect 26065 20893 26099 20927
rect 26433 20893 26467 20927
rect 27445 20893 27479 20927
rect 28917 20893 28951 20927
rect 29009 20893 29043 20927
rect 30674 20893 30708 20927
rect 30941 20893 30975 20927
rect 31217 20893 31251 20927
rect 9413 20825 9447 20859
rect 11069 20825 11103 20859
rect 12909 20825 12943 20859
rect 26249 20825 26283 20859
rect 26341 20825 26375 20859
rect 27353 20825 27387 20859
rect 28181 20825 28215 20859
rect 7389 20757 7423 20791
rect 9321 20757 9355 20791
rect 14197 20757 14231 20791
rect 25329 20757 25363 20791
rect 26985 20757 27019 20791
rect 31033 20757 31067 20791
rect 9229 20553 9263 20587
rect 14657 20553 14691 20587
rect 25053 20553 25087 20587
rect 25513 20553 25547 20587
rect 27905 20553 27939 20587
rect 29285 20553 29319 20587
rect 8493 20485 8527 20519
rect 13185 20485 13219 20519
rect 30420 20485 30454 20519
rect 7481 20417 7515 20451
rect 8677 20417 8711 20451
rect 9505 20417 9539 20451
rect 9597 20417 9631 20451
rect 9689 20417 9723 20451
rect 9873 20417 9907 20451
rect 23673 20417 23707 20451
rect 23940 20417 23974 20451
rect 25605 20417 25639 20451
rect 26525 20417 26559 20451
rect 28457 20417 28491 20451
rect 30665 20417 30699 20451
rect 7665 20349 7699 20383
rect 12909 20349 12943 20383
rect 25697 20349 25731 20383
rect 26985 20349 27019 20383
rect 27261 20349 27295 20383
rect 9321 20281 9355 20315
rect 7297 20213 7331 20247
rect 25145 20213 25179 20247
rect 26341 20213 26375 20247
rect 24041 20009 24075 20043
rect 27445 20009 27479 20043
rect 28549 20009 28583 20043
rect 31401 20009 31435 20043
rect 8401 19941 8435 19975
rect 4445 19873 4479 19907
rect 9505 19873 9539 19907
rect 18981 19873 19015 19907
rect 22017 19873 22051 19907
rect 5457 19805 5491 19839
rect 7021 19805 7055 19839
rect 7288 19805 7322 19839
rect 11989 19805 12023 19839
rect 12265 19805 12299 19839
rect 13369 19805 13403 19839
rect 17693 19805 17727 19839
rect 20729 19805 20763 19839
rect 21189 19805 21223 19839
rect 22845 19805 22879 19839
rect 24225 19805 24259 19839
rect 26065 19805 26099 19839
rect 26332 19805 26366 19839
rect 28728 19805 28762 19839
rect 28825 19805 28859 19839
rect 29100 19805 29134 19839
rect 29193 19805 29227 19839
rect 31217 19805 31251 19839
rect 4169 19737 4203 19771
rect 4813 19737 4847 19771
rect 21833 19737 21867 19771
rect 22293 19737 22327 19771
rect 28917 19737 28951 19771
rect 3801 19669 3835 19703
rect 4261 19669 4295 19703
rect 8953 19669 8987 19703
rect 11345 19669 11379 19703
rect 12081 19669 12115 19703
rect 12817 19669 12851 19703
rect 17509 19669 17543 19703
rect 18337 19669 18371 19703
rect 20177 19669 20211 19703
rect 21005 19669 21039 19703
rect 21465 19669 21499 19703
rect 21925 19669 21959 19703
rect 3893 19465 3927 19499
rect 5365 19465 5399 19499
rect 7849 19465 7883 19499
rect 8217 19465 8251 19499
rect 11345 19465 11379 19499
rect 12909 19465 12943 19499
rect 18613 19465 18647 19499
rect 19257 19465 19291 19499
rect 19625 19465 19659 19499
rect 21649 19465 21683 19499
rect 26985 19465 27019 19499
rect 11796 19397 11830 19431
rect 14933 19397 14967 19431
rect 17500 19397 17534 19431
rect 20536 19397 20570 19431
rect 27261 19397 27295 19431
rect 2513 19329 2547 19363
rect 2780 19329 2814 19363
rect 3985 19329 4019 19363
rect 4252 19329 4286 19363
rect 6009 19329 6043 19363
rect 6377 19329 6411 19363
rect 6633 19329 6667 19363
rect 9965 19329 9999 19363
rect 10232 19329 10266 19363
rect 11529 19329 11563 19363
rect 13369 19329 13403 19363
rect 13829 19329 13863 19363
rect 14841 19329 14875 19363
rect 15117 19329 15151 19363
rect 17233 19329 17267 19363
rect 18889 19329 18923 19363
rect 20269 19329 20303 19363
rect 22946 19329 22980 19363
rect 23213 19329 23247 19363
rect 25973 19329 26007 19363
rect 26433 19329 26467 19363
rect 27164 19329 27198 19363
rect 27353 19329 27387 19363
rect 27536 19329 27570 19363
rect 27629 19329 27663 19363
rect 8309 19261 8343 19295
rect 8401 19261 8435 19295
rect 13461 19261 13495 19295
rect 13645 19261 13679 19295
rect 14381 19261 14415 19295
rect 19717 19261 19751 19295
rect 19901 19261 19935 19295
rect 6193 19193 6227 19227
rect 7757 19193 7791 19227
rect 13001 19125 13035 19159
rect 15301 19125 15335 19159
rect 19073 19125 19107 19159
rect 21833 19125 21867 19159
rect 25789 19125 25823 19159
rect 26617 19125 26651 19159
rect 3065 18921 3099 18955
rect 5917 18921 5951 18955
rect 6653 18921 6687 18955
rect 10609 18921 10643 18955
rect 13185 18921 13219 18955
rect 16129 18921 16163 18955
rect 17601 18921 17635 18955
rect 20637 18921 20671 18955
rect 21189 18921 21223 18955
rect 28365 18921 28399 18955
rect 2973 18853 3007 18887
rect 10885 18853 10919 18887
rect 13921 18853 13955 18887
rect 17141 18853 17175 18887
rect 21097 18853 21131 18887
rect 4445 18785 4479 18819
rect 5181 18785 5215 18819
rect 7113 18785 7147 18819
rect 7297 18785 7331 18819
rect 8033 18785 8067 18819
rect 11437 18785 11471 18819
rect 11805 18785 11839 18819
rect 16773 18785 16807 18819
rect 18245 18785 18279 18819
rect 21649 18785 21683 18819
rect 21833 18785 21867 18819
rect 22569 18785 22603 18819
rect 1409 18717 1443 18751
rect 2789 18717 2823 18751
rect 3249 18717 3283 18751
rect 5365 18717 5399 18751
rect 5641 18717 5675 18751
rect 5733 18717 5767 18751
rect 10793 18717 10827 18751
rect 11253 18717 11287 18751
rect 13277 18717 13311 18751
rect 13370 18717 13404 18751
rect 13783 18717 13817 18751
rect 14473 18717 14507 18751
rect 14749 18717 14783 18751
rect 16957 18717 16991 18751
rect 17969 18717 18003 18751
rect 18521 18717 18555 18751
rect 19257 18717 19291 18751
rect 20913 18717 20947 18751
rect 22937 18717 22971 18751
rect 23305 18717 23339 18751
rect 25513 18717 25547 18751
rect 26985 18717 27019 18751
rect 29009 18717 29043 18751
rect 4169 18649 4203 18683
rect 4629 18649 4663 18683
rect 5549 18649 5583 18683
rect 7021 18649 7055 18683
rect 7481 18649 7515 18683
rect 12050 18649 12084 18683
rect 13553 18649 13587 18683
rect 13645 18649 13679 18683
rect 14994 18649 15028 18683
rect 18061 18649 18095 18683
rect 19502 18649 19536 18683
rect 21557 18649 21591 18683
rect 22017 18649 22051 18683
rect 23029 18649 23063 18683
rect 23121 18649 23155 18683
rect 25780 18649 25814 18683
rect 27230 18649 27264 18683
rect 1593 18581 1627 18615
rect 3801 18581 3835 18615
rect 4261 18581 4295 18615
rect 11345 18581 11379 18615
rect 14657 18581 14691 18615
rect 16221 18581 16255 18615
rect 19073 18581 19107 18615
rect 22753 18581 22787 18615
rect 26893 18581 26927 18615
rect 28457 18581 28491 18615
rect 7849 18377 7883 18411
rect 11897 18377 11931 18411
rect 12173 18377 12207 18411
rect 12541 18377 12575 18411
rect 15117 18377 15151 18411
rect 15485 18377 15519 18411
rect 17233 18377 17267 18411
rect 19165 18377 19199 18411
rect 21649 18377 21683 18411
rect 25973 18377 26007 18411
rect 26341 18377 26375 18411
rect 12633 18309 12667 18343
rect 15577 18309 15611 18343
rect 17570 18309 17604 18343
rect 19257 18309 19291 18343
rect 20085 18309 20119 18343
rect 29193 18309 29227 18343
rect 7665 18241 7699 18275
rect 8217 18241 8251 18275
rect 8677 18241 8711 18275
rect 12081 18241 12115 18275
rect 14298 18241 14332 18275
rect 17049 18241 17083 18275
rect 17325 18241 17359 18275
rect 19993 18241 20027 18275
rect 20453 18241 20487 18275
rect 21189 18241 21223 18275
rect 21465 18241 21499 18275
rect 27353 18241 27387 18275
rect 27905 18241 27939 18275
rect 28457 18241 28491 18275
rect 29653 18241 29687 18275
rect 8309 18173 8343 18207
rect 8493 18173 8527 18207
rect 9229 18173 9263 18207
rect 12817 18173 12851 18207
rect 14565 18173 14599 18207
rect 15669 18173 15703 18207
rect 19349 18173 19383 18207
rect 20269 18173 20303 18207
rect 21005 18173 21039 18207
rect 21281 18173 21315 18207
rect 26433 18173 26467 18207
rect 26617 18173 26651 18207
rect 27445 18173 27479 18207
rect 27537 18173 27571 18207
rect 18797 18105 18831 18139
rect 29377 18105 29411 18139
rect 7481 18037 7515 18071
rect 13185 18037 13219 18071
rect 18705 18037 18739 18071
rect 19625 18037 19659 18071
rect 21465 18037 21499 18071
rect 26985 18037 27019 18071
rect 29745 18037 29779 18071
rect 8401 17833 8435 17867
rect 12725 17833 12759 17867
rect 14289 17833 14323 17867
rect 21005 17833 21039 17867
rect 16313 17765 16347 17799
rect 16405 17765 16439 17799
rect 19809 17765 19843 17799
rect 30665 17765 30699 17799
rect 13277 17697 13311 17731
rect 13461 17697 13495 17731
rect 15025 17697 15059 17731
rect 29377 17697 29411 17731
rect 29745 17697 29779 17731
rect 5641 17629 5675 17663
rect 5825 17629 5859 17663
rect 6193 17629 6227 17663
rect 7021 17629 7055 17663
rect 7288 17629 7322 17663
rect 12173 17629 12207 17663
rect 12449 17629 12483 17663
rect 12541 17629 12575 17663
rect 14105 17629 14139 17663
rect 15853 17629 15887 17663
rect 16037 17629 16071 17663
rect 16221 17629 16255 17663
rect 16497 17629 16531 17663
rect 19257 17629 19291 17663
rect 19441 17629 19475 17663
rect 19533 17629 19567 17663
rect 19625 17629 19659 17663
rect 20453 17629 20487 17663
rect 20729 17629 20763 17663
rect 20821 17629 20855 17663
rect 24409 17629 24443 17663
rect 30849 17629 30883 17663
rect 6009 17561 6043 17595
rect 6101 17561 6135 17595
rect 12357 17561 12391 17595
rect 14841 17561 14875 17595
rect 15301 17561 15335 17595
rect 18429 17561 18463 17595
rect 20637 17561 20671 17595
rect 5089 17493 5123 17527
rect 6377 17493 6411 17527
rect 13553 17493 13587 17527
rect 13921 17493 13955 17527
rect 14473 17493 14507 17527
rect 14933 17493 14967 17527
rect 17141 17493 17175 17527
rect 25053 17493 25087 17527
rect 28733 17493 28767 17527
rect 29837 17493 29871 17527
rect 29929 17493 29963 17527
rect 30297 17493 30331 17527
rect 4813 17289 4847 17323
rect 5273 17289 5307 17323
rect 13277 17289 13311 17323
rect 13369 17289 13403 17323
rect 15485 17289 15519 17323
rect 16313 17289 16347 17323
rect 19073 17289 19107 17323
rect 24869 17289 24903 17323
rect 28457 17289 28491 17323
rect 28917 17289 28951 17323
rect 30389 17289 30423 17323
rect 31125 17289 31159 17323
rect 6828 17221 6862 17255
rect 8861 17221 8895 17255
rect 14350 17221 14384 17255
rect 15945 17221 15979 17255
rect 16129 17221 16163 17255
rect 28365 17221 28399 17255
rect 30052 17221 30086 17255
rect 3433 17153 3467 17187
rect 3689 17153 3723 17187
rect 8769 17153 8803 17187
rect 9045 17153 9079 17187
rect 10425 17153 10459 17187
rect 13093 17153 13127 17187
rect 14105 17153 14139 17187
rect 17693 17153 17727 17187
rect 17960 17153 17994 17187
rect 22477 17153 22511 17187
rect 23857 17153 23891 17187
rect 24777 17153 24811 17187
rect 26249 17153 26283 17187
rect 26341 17153 26375 17187
rect 26433 17153 26467 17187
rect 26617 17153 26651 17187
rect 30297 17153 30331 17187
rect 31309 17153 31343 17187
rect 5365 17085 5399 17119
rect 5457 17085 5491 17119
rect 6561 17085 6595 17119
rect 8677 17085 8711 17119
rect 13921 17085 13955 17119
rect 23581 17085 23615 17119
rect 24593 17085 24627 17119
rect 25881 17085 25915 17119
rect 28273 17085 28307 17119
rect 30941 17085 30975 17119
rect 7941 17017 7975 17051
rect 25237 17017 25271 17051
rect 4905 16949 4939 16983
rect 8033 16949 8067 16983
rect 9229 16949 9263 16983
rect 10241 16949 10275 16983
rect 22293 16949 22327 16983
rect 22937 16949 22971 16983
rect 24041 16949 24075 16983
rect 25329 16949 25363 16983
rect 26065 16949 26099 16983
rect 28825 16949 28859 16983
rect 3341 16745 3375 16779
rect 6929 16745 6963 16779
rect 18245 16745 18279 16779
rect 24225 16745 24259 16779
rect 25789 16745 25823 16779
rect 11161 16677 11195 16711
rect 28733 16677 28767 16711
rect 3801 16609 3835 16643
rect 5917 16609 5951 16643
rect 7757 16609 7791 16643
rect 9781 16609 9815 16643
rect 11805 16609 11839 16643
rect 23581 16609 23615 16643
rect 24409 16609 24443 16643
rect 29561 16609 29595 16643
rect 3157 16541 3191 16575
rect 3433 16541 3467 16575
rect 7113 16541 7147 16575
rect 7573 16541 7607 16575
rect 10048 16541 10082 16575
rect 18429 16541 18463 16575
rect 21833 16541 21867 16575
rect 22100 16541 22134 16575
rect 23765 16541 23799 16575
rect 26065 16541 26099 16575
rect 28912 16541 28946 16575
rect 29009 16541 29043 16575
rect 29284 16541 29318 16575
rect 29377 16541 29411 16575
rect 29828 16541 29862 16575
rect 4046 16473 4080 16507
rect 5273 16473 5307 16507
rect 7665 16473 7699 16507
rect 24654 16473 24688 16507
rect 29101 16473 29135 16507
rect 3617 16405 3651 16439
rect 5181 16405 5215 16439
rect 7205 16405 7239 16439
rect 11253 16405 11287 16439
rect 23213 16405 23247 16439
rect 23857 16405 23891 16439
rect 25881 16405 25915 16439
rect 30941 16405 30975 16439
rect 4261 16201 4295 16235
rect 4629 16201 4663 16235
rect 4721 16201 4755 16235
rect 10517 16201 10551 16235
rect 10885 16201 10919 16235
rect 21649 16201 21683 16235
rect 23857 16201 23891 16235
rect 27261 16201 27295 16235
rect 9229 16133 9263 16167
rect 11529 16133 11563 16167
rect 11713 16133 11747 16167
rect 22078 16133 22112 16167
rect 23489 16133 23523 16167
rect 23581 16133 23615 16167
rect 25084 16133 25118 16167
rect 25973 16133 26007 16167
rect 8953 16065 8987 16099
rect 9046 16065 9080 16099
rect 9321 16065 9355 16099
rect 9459 16065 9493 16099
rect 9965 16065 9999 16099
rect 10241 16065 10275 16099
rect 11897 16065 11931 16099
rect 15209 16065 15243 16099
rect 21465 16065 21499 16099
rect 23305 16065 23339 16099
rect 23673 16065 23707 16099
rect 25697 16065 25731 16099
rect 25789 16065 25823 16099
rect 26341 16065 26375 16099
rect 27353 16065 27387 16099
rect 27813 16065 27847 16099
rect 4813 15997 4847 16031
rect 10149 15997 10183 16031
rect 10977 15997 11011 16031
rect 11069 15997 11103 16031
rect 21833 15997 21867 16031
rect 25329 15997 25363 16031
rect 27077 15997 27111 16031
rect 28365 15997 28399 16031
rect 9597 15929 9631 15963
rect 10057 15929 10091 15963
rect 23213 15929 23247 15963
rect 25513 15929 25547 15963
rect 10425 15861 10459 15895
rect 15485 15861 15519 15895
rect 23949 15861 23983 15895
rect 25973 15861 26007 15895
rect 26525 15861 26559 15895
rect 27721 15861 27755 15895
rect 8309 15657 8343 15691
rect 10333 15657 10367 15691
rect 22477 15657 22511 15691
rect 26157 15657 26191 15691
rect 8769 15589 8803 15623
rect 8953 15521 8987 15555
rect 10977 15521 11011 15555
rect 22937 15521 22971 15555
rect 23029 15521 23063 15555
rect 23857 15521 23891 15555
rect 25513 15521 25547 15555
rect 7205 15453 7239 15487
rect 7757 15453 7791 15487
rect 8033 15453 8067 15487
rect 8125 15453 8159 15487
rect 8585 15453 8619 15487
rect 10425 15453 10459 15487
rect 11989 15453 12023 15487
rect 12633 15453 12667 15487
rect 17785 15453 17819 15487
rect 18153 15453 18187 15487
rect 18429 15453 18463 15487
rect 19901 15453 19935 15487
rect 20453 15453 20487 15487
rect 20637 15453 20671 15487
rect 20821 15453 20855 15487
rect 26249 15453 26283 15487
rect 28273 15453 28307 15487
rect 28641 15453 28675 15487
rect 7941 15385 7975 15419
rect 9198 15385 9232 15419
rect 19257 15385 19291 15419
rect 20729 15385 20763 15419
rect 22845 15385 22879 15419
rect 23305 15385 23339 15419
rect 25697 15385 25731 15419
rect 26516 15385 26550 15419
rect 27721 15385 27755 15419
rect 6653 15317 6687 15351
rect 17601 15317 17635 15351
rect 18337 15317 18371 15351
rect 18613 15317 18647 15351
rect 21005 15317 21039 15351
rect 25789 15317 25823 15351
rect 27629 15317 27663 15351
rect 28457 15317 28491 15351
rect 3065 15113 3099 15147
rect 6745 15113 6779 15147
rect 6837 15113 6871 15147
rect 8033 15113 8067 15147
rect 8861 15113 8895 15147
rect 9229 15113 9263 15147
rect 22201 15113 22235 15147
rect 22569 15113 22603 15147
rect 26249 15113 26283 15147
rect 26985 15113 27019 15147
rect 9321 15045 9355 15079
rect 12440 15045 12474 15079
rect 26525 15045 26559 15079
rect 2881 14977 2915 15011
rect 3433 14977 3467 15011
rect 3893 14977 3927 15011
rect 7941 14977 7975 15011
rect 14933 14977 14967 15011
rect 17325 14977 17359 15011
rect 17592 14977 17626 15011
rect 18797 14977 18831 15011
rect 19053 14977 19087 15011
rect 22017 14977 22051 15011
rect 22661 14977 22695 15011
rect 26433 14977 26467 15011
rect 26617 14977 26651 15011
rect 26801 14977 26835 15011
rect 28109 14977 28143 15011
rect 28365 14977 28399 15011
rect 3525 14909 3559 14943
rect 3709 14909 3743 14943
rect 4537 14909 4571 14943
rect 7021 14909 7055 14943
rect 8217 14909 8251 14943
rect 9505 14909 9539 14943
rect 12173 14909 12207 14943
rect 14197 14909 14231 14943
rect 20821 14909 20855 14943
rect 21005 14909 21039 14943
rect 22753 14909 22787 14943
rect 20177 14841 20211 14875
rect 21833 14841 21867 14875
rect 2697 14773 2731 14807
rect 6377 14773 6411 14807
rect 7573 14773 7607 14807
rect 13553 14773 13587 14807
rect 13645 14773 13679 14807
rect 14381 14773 14415 14807
rect 18705 14773 18739 14807
rect 20269 14773 20303 14807
rect 21649 14773 21683 14807
rect 6377 14569 6411 14603
rect 7849 14569 7883 14603
rect 7941 14569 7975 14603
rect 12449 14569 12483 14603
rect 17877 14569 17911 14603
rect 19257 14569 19291 14603
rect 12725 14501 12759 14535
rect 16037 14501 16071 14535
rect 4445 14433 4479 14467
rect 10609 14433 10643 14467
rect 13369 14433 13403 14467
rect 14657 14433 14691 14467
rect 16681 14433 16715 14467
rect 17233 14433 17267 14467
rect 18337 14433 18371 14467
rect 18521 14433 18555 14467
rect 19901 14433 19935 14467
rect 2237 14365 2271 14399
rect 4997 14365 5031 14399
rect 6469 14365 6503 14399
rect 8493 14365 8527 14399
rect 12633 14365 12667 14399
rect 13093 14365 13127 14399
rect 13737 14365 13771 14399
rect 14381 14365 14415 14399
rect 17417 14365 17451 14399
rect 19625 14365 19659 14399
rect 21382 14365 21416 14399
rect 21649 14365 21683 14399
rect 2504 14297 2538 14331
rect 5264 14297 5298 14331
rect 6736 14297 6770 14331
rect 10876 14297 10910 14331
rect 13185 14297 13219 14331
rect 14902 14297 14936 14331
rect 19717 14297 19751 14331
rect 3617 14229 3651 14263
rect 3801 14229 3835 14263
rect 4169 14229 4203 14263
rect 4261 14229 4295 14263
rect 11989 14229 12023 14263
rect 13553 14229 13587 14263
rect 14565 14229 14599 14263
rect 16129 14229 16163 14263
rect 17325 14229 17359 14263
rect 17785 14229 17819 14263
rect 18245 14229 18279 14263
rect 20269 14229 20303 14263
rect 3709 14025 3743 14059
rect 3985 14025 4019 14059
rect 6009 14025 6043 14059
rect 7021 14025 7055 14059
rect 10977 14025 11011 14059
rect 11529 14025 11563 14059
rect 11897 14025 11931 14059
rect 12449 14025 12483 14059
rect 13921 14025 13955 14059
rect 14289 14025 14323 14059
rect 14933 14025 14967 14059
rect 15301 14025 15335 14059
rect 19717 14025 19751 14059
rect 20361 14025 20395 14059
rect 21097 14025 21131 14059
rect 22293 14025 22327 14059
rect 2596 13957 2630 13991
rect 4997 13957 5031 13991
rect 13562 13957 13596 13991
rect 15945 13957 15979 13991
rect 18604 13957 18638 13991
rect 19993 13957 20027 13991
rect 20085 13957 20119 13991
rect 25053 13957 25087 13991
rect 2329 13889 2363 13923
rect 4537 13889 4571 13923
rect 4721 13889 4755 13923
rect 4905 13889 4939 13923
rect 5089 13889 5123 13923
rect 6193 13889 6227 13923
rect 7205 13889 7239 13923
rect 11161 13889 11195 13923
rect 15761 13889 15795 13923
rect 16681 13889 16715 13923
rect 18337 13889 18371 13923
rect 19809 13889 19843 13923
rect 20177 13889 20211 13923
rect 21005 13889 21039 13923
rect 21833 13889 21867 13923
rect 22017 13889 22051 13923
rect 22109 13889 22143 13923
rect 24961 13889 24995 13923
rect 25145 13889 25179 13923
rect 25329 13889 25363 13923
rect 25973 13889 26007 13923
rect 26341 13889 26375 13923
rect 27905 13889 27939 13923
rect 29009 13889 29043 13923
rect 29469 13889 29503 13923
rect 31217 13889 31251 13923
rect 11989 13821 12023 13855
rect 12081 13821 12115 13855
rect 13829 13821 13863 13855
rect 14381 13821 14415 13855
rect 14473 13821 14507 13855
rect 15393 13821 15427 13855
rect 15577 13821 15611 13855
rect 20821 13821 20855 13855
rect 29101 13821 29135 13855
rect 29285 13821 29319 13855
rect 30113 13821 30147 13855
rect 31493 13821 31527 13855
rect 5273 13753 5307 13787
rect 16865 13753 16899 13787
rect 21465 13753 21499 13787
rect 24777 13753 24811 13787
rect 16129 13685 16163 13719
rect 22017 13685 22051 13719
rect 25421 13685 25455 13719
rect 26157 13685 26191 13719
rect 27353 13685 27387 13719
rect 28641 13685 28675 13719
rect 3801 13481 3835 13515
rect 14105 13481 14139 13515
rect 19257 13481 19291 13515
rect 25789 13481 25823 13515
rect 27261 13481 27295 13515
rect 29377 13481 29411 13515
rect 13921 13413 13955 13447
rect 14565 13345 14599 13379
rect 14657 13345 14691 13379
rect 15485 13345 15519 13379
rect 19809 13345 19843 13379
rect 3985 13277 4019 13311
rect 12265 13277 12299 13311
rect 12541 13277 12575 13311
rect 15853 13277 15887 13311
rect 15945 13277 15979 13311
rect 16037 13277 16071 13311
rect 16129 13277 16163 13311
rect 16313 13277 16347 13311
rect 16589 13277 16623 13311
rect 24041 13277 24075 13311
rect 24409 13277 24443 13311
rect 25881 13277 25915 13311
rect 27721 13277 27755 13311
rect 27997 13277 28031 13311
rect 29699 13277 29733 13311
rect 30112 13277 30146 13311
rect 30205 13277 30239 13311
rect 12786 13209 12820 13243
rect 14473 13209 14507 13243
rect 14933 13209 14967 13243
rect 16773 13209 16807 13243
rect 24654 13209 24688 13243
rect 26148 13209 26182 13243
rect 28242 13209 28276 13243
rect 29837 13209 29871 13243
rect 29929 13209 29963 13243
rect 12449 13141 12483 13175
rect 15669 13141 15703 13175
rect 16405 13141 16439 13175
rect 24225 13141 24259 13175
rect 27905 13141 27939 13175
rect 29561 13141 29595 13175
rect 10425 12937 10459 12971
rect 14289 12937 14323 12971
rect 24501 12937 24535 12971
rect 24869 12937 24903 12971
rect 26985 12937 27019 12971
rect 27353 12937 27387 12971
rect 28549 12937 28583 12971
rect 30021 12937 30055 12971
rect 1777 12869 1811 12903
rect 10609 12869 10643 12903
rect 13001 12869 13035 12903
rect 13921 12869 13955 12903
rect 24961 12869 24995 12903
rect 26709 12869 26743 12903
rect 28886 12869 28920 12903
rect 8677 12801 8711 12835
rect 10701 12801 10735 12835
rect 12817 12801 12851 12835
rect 13093 12801 13127 12835
rect 13185 12801 13219 12835
rect 13645 12801 13679 12835
rect 13738 12801 13772 12835
rect 14013 12801 14047 12835
rect 14151 12801 14185 12835
rect 20545 12801 20579 12835
rect 22201 12801 22235 12835
rect 25881 12801 25915 12835
rect 27445 12801 27479 12835
rect 28365 12801 28399 12835
rect 28641 12801 28675 12835
rect 30665 12801 30699 12835
rect 8953 12733 8987 12767
rect 21373 12733 21407 12767
rect 23857 12733 23891 12767
rect 25145 12733 25179 12767
rect 27537 12733 27571 12767
rect 13369 12665 13403 12699
rect 1501 12597 1535 12631
rect 22017 12597 22051 12631
rect 23305 12597 23339 12631
rect 30113 12597 30147 12631
rect 9137 12393 9171 12427
rect 22937 12393 22971 12427
rect 29561 12393 29595 12427
rect 6101 12257 6135 12291
rect 6285 12257 6319 12291
rect 9965 12257 9999 12291
rect 15669 12257 15703 12291
rect 15853 12257 15887 12291
rect 19901 12257 19935 12291
rect 21465 12257 21499 12291
rect 23581 12257 23615 12291
rect 30021 12257 30055 12291
rect 30205 12257 30239 12291
rect 4905 12189 4939 12223
rect 5181 12189 5215 12223
rect 7021 12189 7055 12223
rect 8033 12189 8067 12223
rect 8677 12189 8711 12223
rect 9321 12189 9355 12223
rect 9781 12189 9815 12223
rect 16957 12189 16991 12223
rect 20821 12189 20855 12223
rect 21189 12189 21223 12223
rect 23305 12189 23339 12223
rect 15945 12121 15979 12155
rect 16405 12121 16439 12155
rect 19625 12121 19659 12155
rect 20177 12121 20211 12155
rect 21710 12121 21744 12155
rect 25421 12121 25455 12155
rect 26157 12121 26191 12155
rect 29929 12121 29963 12155
rect 4261 12053 4295 12087
rect 4997 12053 5031 12087
rect 6377 12053 6411 12087
rect 6745 12053 6779 12087
rect 6837 12053 6871 12087
rect 7389 12053 7423 12087
rect 8493 12053 8527 12087
rect 9413 12053 9447 12087
rect 9873 12053 9907 12087
rect 16313 12053 16347 12087
rect 19257 12053 19291 12087
rect 19717 12053 19751 12087
rect 21373 12053 21407 12087
rect 22845 12053 22879 12087
rect 23397 12053 23431 12087
rect 3985 11849 4019 11883
rect 4445 11849 4479 11883
rect 4813 11849 4847 11883
rect 6193 11849 6227 11883
rect 7757 11849 7791 11883
rect 16497 11849 16531 11883
rect 23213 11849 23247 11883
rect 6644 11781 6678 11815
rect 8125 11781 8159 11815
rect 21557 11781 21591 11815
rect 22100 11781 22134 11815
rect 23305 11781 23339 11815
rect 26525 11781 26559 11815
rect 2605 11713 2639 11747
rect 2872 11713 2906 11747
rect 4905 11713 4939 11747
rect 5089 11713 5123 11747
rect 5181 11713 5215 11747
rect 5273 11713 5307 11747
rect 6377 11713 6411 11747
rect 7849 11713 7883 11747
rect 8033 11713 8067 11747
rect 8217 11713 8251 11747
rect 9413 11713 9447 11747
rect 13737 11713 13771 11747
rect 15384 11713 15418 11747
rect 17960 11713 17994 11747
rect 19432 11713 19466 11747
rect 20821 11713 20855 11747
rect 21833 11713 21867 11747
rect 23857 11713 23891 11747
rect 25789 11713 25823 11747
rect 26341 11713 26375 11747
rect 26433 11713 26467 11747
rect 26709 11713 26743 11747
rect 27537 11713 27571 11747
rect 4169 11645 4203 11679
rect 4353 11645 4387 11679
rect 5641 11645 5675 11679
rect 8677 11645 8711 11679
rect 15117 11645 15151 11679
rect 17693 11645 17727 11679
rect 19165 11645 19199 11679
rect 5457 11509 5491 11543
rect 8401 11509 8435 11543
rect 13921 11509 13955 11543
rect 19073 11509 19107 11543
rect 20545 11509 20579 11543
rect 25605 11509 25639 11543
rect 26157 11509 26191 11543
rect 26985 11509 27019 11543
rect 5549 11305 5583 11339
rect 18061 11305 18095 11339
rect 18797 11305 18831 11339
rect 21925 11305 21959 11339
rect 22753 11305 22787 11339
rect 26617 11305 26651 11339
rect 28089 11305 28123 11339
rect 2145 11237 2179 11271
rect 3801 11237 3835 11271
rect 8769 11237 8803 11271
rect 16313 11237 16347 11271
rect 19257 11237 19291 11271
rect 2237 11169 2271 11203
rect 4261 11169 4295 11203
rect 4353 11169 4387 11203
rect 7389 11169 7423 11203
rect 10517 11169 10551 11203
rect 11713 11169 11747 11203
rect 19901 11169 19935 11203
rect 20729 11169 20763 11203
rect 22569 11169 22603 11203
rect 28733 11169 28767 11203
rect 1961 11101 1995 11135
rect 2493 11101 2527 11135
rect 5181 11101 5215 11135
rect 6929 11101 6963 11135
rect 7205 11101 7239 11135
rect 9045 11101 9079 11135
rect 10885 11101 10919 11135
rect 13001 11101 13035 11135
rect 14105 11101 14139 11135
rect 14361 11101 14395 11135
rect 16129 11101 16163 11135
rect 16497 11101 16531 11135
rect 18245 11101 18279 11135
rect 18613 11101 18647 11135
rect 21005 11101 21039 11135
rect 21373 11101 21407 11135
rect 22293 11101 22327 11135
rect 22937 11101 22971 11135
rect 23029 11101 23063 11135
rect 23305 11101 23339 11135
rect 25237 11101 25271 11135
rect 26709 11101 26743 11135
rect 4169 11033 4203 11067
rect 4629 11033 4663 11067
rect 6684 11033 6718 11067
rect 7656 11033 7690 11067
rect 9873 11033 9907 11067
rect 13737 11033 13771 11067
rect 19625 11033 19659 11067
rect 20085 11033 20119 11067
rect 21097 11033 21131 11067
rect 21189 11033 21223 11067
rect 23121 11033 23155 11067
rect 25504 11033 25538 11067
rect 26954 11033 26988 11067
rect 3617 10965 3651 10999
rect 7021 10965 7055 10999
rect 9965 10965 9999 10999
rect 10701 10965 10735 10999
rect 12357 10965 12391 10999
rect 15485 10965 15519 10999
rect 15577 10965 15611 10999
rect 19717 10965 19751 10999
rect 20821 10965 20855 10999
rect 22385 10965 22419 10999
rect 28181 10965 28215 10999
rect 6101 10761 6135 10795
rect 6929 10761 6963 10795
rect 7297 10761 7331 10795
rect 8217 10761 8251 10795
rect 8493 10761 8527 10795
rect 8953 10761 8987 10795
rect 9321 10761 9355 10795
rect 11345 10761 11379 10795
rect 11529 10761 11563 10795
rect 11897 10761 11931 10795
rect 14197 10761 14231 10795
rect 14565 10761 14599 10795
rect 25697 10761 25731 10795
rect 26065 10761 26099 10795
rect 26709 10761 26743 10795
rect 27353 10761 27387 10795
rect 4445 10693 4479 10727
rect 5825 10693 5859 10727
rect 6837 10693 6871 10727
rect 10232 10693 10266 10727
rect 13001 10693 13035 10727
rect 13829 10693 13863 10727
rect 2769 10625 2803 10659
rect 4353 10625 4387 10659
rect 4813 10625 4847 10659
rect 5549 10625 5583 10659
rect 5733 10625 5767 10659
rect 5917 10625 5951 10659
rect 8033 10625 8067 10659
rect 8309 10625 8343 10659
rect 8401 10625 8435 10659
rect 8677 10625 8711 10659
rect 9413 10625 9447 10659
rect 11989 10625 12023 10659
rect 14657 10625 14691 10659
rect 19625 10625 19659 10659
rect 19901 10625 19935 10659
rect 20361 10625 20395 10659
rect 26525 10625 26559 10659
rect 2513 10557 2547 10591
rect 4629 10557 4663 10591
rect 5365 10557 5399 10591
rect 6653 10557 6687 10591
rect 9505 10557 9539 10591
rect 9965 10557 9999 10591
rect 12173 10557 12207 10591
rect 14841 10557 14875 10591
rect 19717 10557 19751 10591
rect 26157 10557 26191 10591
rect 26249 10557 26283 10591
rect 27445 10557 27479 10591
rect 27537 10557 27571 10591
rect 29929 10557 29963 10591
rect 3893 10489 3927 10523
rect 26985 10489 27019 10523
rect 3985 10421 4019 10455
rect 7849 10421 7883 10455
rect 8861 10421 8895 10455
rect 19901 10421 19935 10455
rect 20085 10421 20119 10455
rect 20177 10421 20211 10455
rect 29285 10421 29319 10455
rect 2605 10217 2639 10251
rect 9965 10217 9999 10251
rect 20913 10217 20947 10251
rect 10241 10149 10275 10183
rect 23857 10149 23891 10183
rect 29561 10149 29595 10183
rect 4353 10081 4387 10115
rect 8493 10081 8527 10115
rect 19993 10081 20027 10115
rect 24961 10081 24995 10115
rect 30113 10081 30147 10115
rect 2789 10013 2823 10047
rect 5181 10013 5215 10047
rect 9505 10013 9539 10047
rect 10149 10013 10183 10047
rect 10333 10013 10367 10047
rect 10425 10013 10459 10047
rect 10793 10013 10827 10047
rect 10977 10013 11011 10047
rect 11713 10013 11747 10047
rect 14105 10013 14139 10047
rect 14381 10013 14415 10047
rect 14841 10013 14875 10047
rect 20729 10013 20763 10047
rect 21092 10013 21126 10047
rect 21409 10013 21443 10047
rect 21557 10013 21591 10047
rect 23673 10013 23707 10047
rect 25881 10013 25915 10047
rect 29101 10013 29135 10047
rect 30389 10013 30423 10047
rect 30482 10013 30516 10047
rect 30854 10013 30888 10047
rect 4169 9945 4203 9979
rect 4629 9945 4663 9979
rect 8309 9945 8343 9979
rect 8953 9945 8987 9979
rect 11161 9945 11195 9979
rect 11897 9945 11931 9979
rect 14197 9945 14231 9979
rect 14565 9945 14599 9979
rect 19717 9945 19751 9979
rect 20177 9945 20211 9979
rect 21189 9945 21223 9979
rect 21281 9945 21315 9979
rect 24777 9945 24811 9979
rect 25237 9945 25271 9979
rect 29929 9945 29963 9979
rect 30665 9945 30699 9979
rect 30757 9945 30791 9979
rect 3801 9877 3835 9911
rect 4261 9877 4295 9911
rect 7941 9877 7975 9911
rect 8401 9877 8435 9911
rect 11529 9877 11563 9911
rect 14657 9877 14691 9911
rect 19349 9877 19383 9911
rect 19809 9877 19843 9911
rect 24409 9877 24443 9911
rect 24869 9877 24903 9911
rect 29285 9877 29319 9911
rect 30021 9877 30055 9911
rect 31033 9877 31067 9911
rect 8401 9673 8435 9707
rect 11345 9673 11379 9707
rect 12909 9673 12943 9707
rect 18797 9673 18831 9707
rect 20269 9673 20303 9707
rect 20361 9673 20395 9707
rect 30205 9673 30239 9707
rect 30481 9673 30515 9707
rect 11774 9605 11808 9639
rect 14188 9605 14222 9639
rect 16129 9605 16163 9639
rect 19134 9605 19168 9639
rect 20821 9605 20855 9639
rect 25114 9605 25148 9639
rect 28273 9605 28307 9639
rect 28365 9605 28399 9639
rect 29092 9605 29126 9639
rect 2513 9537 2547 9571
rect 2780 9537 2814 9571
rect 7288 9537 7322 9571
rect 11161 9537 11195 9571
rect 11529 9537 11563 9571
rect 13553 9537 13587 9571
rect 13921 9537 13955 9571
rect 16313 9537 16347 9571
rect 18613 9537 18647 9571
rect 18889 9537 18923 9571
rect 20729 9537 20763 9571
rect 23121 9537 23155 9571
rect 23397 9537 23431 9571
rect 23653 9537 23687 9571
rect 24869 9537 24903 9571
rect 31033 9537 31067 9571
rect 7021 9469 7055 9503
rect 15945 9469 15979 9503
rect 21005 9469 21039 9503
rect 28181 9469 28215 9503
rect 28832 9469 28866 9503
rect 3893 9401 3927 9435
rect 15301 9401 15335 9435
rect 23305 9401 23339 9435
rect 13001 9333 13035 9367
rect 15393 9333 15427 9367
rect 16497 9333 16531 9367
rect 24777 9333 24811 9367
rect 26249 9333 26283 9367
rect 28733 9333 28767 9367
rect 2881 9129 2915 9163
rect 7481 9129 7515 9163
rect 11897 9129 11931 9163
rect 15117 9129 15151 9163
rect 19073 9129 19107 9163
rect 20821 9129 20855 9163
rect 22845 9129 22879 9163
rect 24409 9129 24443 9163
rect 26433 9129 26467 9163
rect 29193 9129 29227 9163
rect 30941 9129 30975 9163
rect 11253 9061 11287 9095
rect 23029 9061 23063 9095
rect 11161 8993 11195 9027
rect 12541 8993 12575 9027
rect 14565 8993 14599 9027
rect 17601 8993 17635 9027
rect 21373 8993 21407 9027
rect 25053 8993 25087 9027
rect 25789 8993 25823 9027
rect 29561 8993 29595 9027
rect 3065 8925 3099 8959
rect 7665 8925 7699 8959
rect 10149 8925 10183 8959
rect 11069 8925 11103 8959
rect 11345 8925 11379 8959
rect 12265 8925 12299 8959
rect 14749 8925 14783 8959
rect 18337 8925 18371 8959
rect 18521 8925 18555 8959
rect 18797 8925 18831 8959
rect 18889 8925 18923 8959
rect 19349 8925 19383 8959
rect 22753 8925 22787 8959
rect 22845 8925 22879 8959
rect 23760 8925 23794 8959
rect 23857 8925 23891 8959
rect 24132 8925 24166 8959
rect 24225 8925 24259 8959
rect 26617 8925 26651 8959
rect 26709 8925 26743 8959
rect 29009 8925 29043 8959
rect 29817 8925 29851 8959
rect 10885 8857 10919 8891
rect 17325 8857 17359 8891
rect 17785 8857 17819 8891
rect 18705 8857 18739 8891
rect 19616 8857 19650 8891
rect 22569 8857 22603 8891
rect 23949 8857 23983 8891
rect 24777 8857 24811 8891
rect 25237 8857 25271 8891
rect 26433 8857 26467 8891
rect 10793 8789 10827 8823
rect 12357 8789 12391 8823
rect 14657 8789 14691 8823
rect 16957 8789 16991 8823
rect 17417 8789 17451 8823
rect 20729 8789 20763 8823
rect 23581 8789 23615 8823
rect 24869 8789 24903 8823
rect 26893 8789 26927 8823
rect 9873 8585 9907 8619
rect 10517 8585 10551 8619
rect 18061 8585 18095 8619
rect 18153 8585 18187 8619
rect 22477 8585 22511 8619
rect 26249 8585 26283 8619
rect 9597 8517 9631 8551
rect 14197 8517 14231 8551
rect 14289 8517 14323 8551
rect 22109 8517 22143 8551
rect 6009 8449 6043 8483
rect 8125 8449 8159 8483
rect 8309 8449 8343 8483
rect 8401 8449 8435 8483
rect 8493 8449 8527 8483
rect 9229 8449 9263 8483
rect 9322 8449 9356 8483
rect 9505 8449 9539 8483
rect 9735 8449 9769 8483
rect 13921 8449 13955 8483
rect 14069 8449 14103 8483
rect 14386 8449 14420 8483
rect 14657 8449 14691 8483
rect 14841 8449 14875 8483
rect 14933 8449 14967 8483
rect 15117 8449 15151 8483
rect 16037 8449 16071 8483
rect 16313 8449 16347 8483
rect 16681 8449 16715 8483
rect 16937 8449 16971 8483
rect 18521 8449 18555 8483
rect 18981 8449 19015 8483
rect 21925 8449 21959 8483
rect 22201 8449 22235 8483
rect 22293 8449 22327 8483
rect 26433 8449 26467 8483
rect 26525 8449 26559 8483
rect 26617 8449 26651 8483
rect 26801 8449 26835 8483
rect 27445 8449 27479 8483
rect 27905 8449 27939 8483
rect 28457 8449 28491 8483
rect 28641 8449 28675 8483
rect 7389 8381 7423 8415
rect 10609 8381 10643 8415
rect 10793 8381 10827 8415
rect 15025 8381 15059 8415
rect 18613 8381 18647 8415
rect 18797 8381 18831 8415
rect 19533 8381 19567 8415
rect 27169 8381 27203 8415
rect 27353 8381 27387 8415
rect 5825 8313 5859 8347
rect 10149 8313 10183 8347
rect 14565 8313 14599 8347
rect 16221 8313 16255 8347
rect 16497 8313 16531 8347
rect 28825 8313 28859 8347
rect 6837 8245 6871 8279
rect 8677 8245 8711 8279
rect 27813 8245 27847 8279
rect 9781 8041 9815 8075
rect 17969 8041 18003 8075
rect 27537 8041 27571 8075
rect 31125 8041 31159 8075
rect 6653 7973 6687 8007
rect 5273 7905 5307 7939
rect 7389 7905 7423 7939
rect 8125 7905 8159 7939
rect 11161 7905 11195 7939
rect 14657 7905 14691 7939
rect 20637 7905 20671 7939
rect 21557 7905 21591 7939
rect 22569 7905 22603 7939
rect 23397 7905 23431 7939
rect 9045 7837 9079 7871
rect 9138 7837 9172 7871
rect 9321 7837 9355 7871
rect 9413 7837 9447 7871
rect 9551 7837 9585 7871
rect 13553 7837 13587 7871
rect 15485 7837 15519 7871
rect 16589 7837 16623 7871
rect 16856 7837 16890 7871
rect 22385 7837 22419 7871
rect 25789 7837 25823 7871
rect 26065 7837 26099 7871
rect 28917 7837 28951 7871
rect 5540 7769 5574 7803
rect 7113 7769 7147 7803
rect 7573 7769 7607 7803
rect 10894 7769 10928 7803
rect 14473 7769 14507 7803
rect 14933 7769 14967 7803
rect 20453 7769 20487 7803
rect 20913 7769 20947 7803
rect 22293 7769 22327 7803
rect 22845 7769 22879 7803
rect 26310 7769 26344 7803
rect 28650 7769 28684 7803
rect 31401 7769 31435 7803
rect 6745 7701 6779 7735
rect 7205 7701 7239 7735
rect 9689 7701 9723 7735
rect 13369 7701 13403 7735
rect 14105 7701 14139 7735
rect 14565 7701 14599 7735
rect 20085 7701 20119 7735
rect 20545 7701 20579 7735
rect 21925 7701 21959 7735
rect 25973 7701 26007 7735
rect 27445 7701 27479 7735
rect 5641 7497 5675 7531
rect 6377 7497 6411 7531
rect 6745 7497 6779 7531
rect 6837 7497 6871 7531
rect 7665 7497 7699 7531
rect 10425 7497 10459 7531
rect 14565 7497 14599 7531
rect 21649 7497 21683 7531
rect 23213 7497 23247 7531
rect 26985 7497 27019 7531
rect 28733 7497 28767 7531
rect 22078 7429 22112 7463
rect 27445 7429 27479 7463
rect 5825 7361 5859 7395
rect 7573 7361 7607 7395
rect 8033 7361 8067 7395
rect 8769 7361 8803 7395
rect 9034 7361 9068 7395
rect 9301 7361 9335 7395
rect 11069 7361 11103 7395
rect 13441 7361 13475 7395
rect 15025 7361 15059 7395
rect 15485 7361 15519 7395
rect 19533 7361 19567 7395
rect 19809 7361 19843 7395
rect 20065 7361 20099 7395
rect 21465 7361 21499 7395
rect 21833 7361 21867 7395
rect 27353 7361 27387 7395
rect 28549 7361 28583 7395
rect 7021 7293 7055 7327
rect 7849 7293 7883 7327
rect 8585 7293 8619 7327
rect 13185 7293 13219 7327
rect 15117 7293 15151 7327
rect 15209 7293 15243 7327
rect 16037 7293 16071 7327
rect 27537 7293 27571 7327
rect 27813 7293 27847 7327
rect 28365 7293 28399 7327
rect 8953 7225 8987 7259
rect 19717 7225 19751 7259
rect 7205 7157 7239 7191
rect 10517 7157 10551 7191
rect 14657 7157 14691 7191
rect 21189 7157 21223 7191
rect 9505 6953 9539 6987
rect 10701 6953 10735 6987
rect 15485 6953 15519 6987
rect 13737 6885 13771 6919
rect 5457 6817 5491 6851
rect 10057 6817 10091 6851
rect 24961 6817 24995 6851
rect 6929 6749 6963 6783
rect 10517 6749 10551 6783
rect 13185 6749 13219 6783
rect 13553 6749 13587 6783
rect 14105 6749 14139 6783
rect 17141 6749 17175 6783
rect 23949 6749 23983 6783
rect 25789 6749 25823 6783
rect 25973 6749 26007 6783
rect 26341 6749 26375 6783
rect 5724 6681 5758 6715
rect 7174 6681 7208 6715
rect 9965 6681 9999 6715
rect 13369 6681 13403 6715
rect 13461 6681 13495 6715
rect 14350 6681 14384 6715
rect 16681 6681 16715 6715
rect 24777 6681 24811 6715
rect 25237 6681 25271 6715
rect 26157 6681 26191 6715
rect 26249 6681 26283 6715
rect 6837 6613 6871 6647
rect 8309 6613 8343 6647
rect 9873 6613 9907 6647
rect 16773 6613 16807 6647
rect 17325 6613 17359 6647
rect 24133 6613 24167 6647
rect 24409 6613 24443 6647
rect 24869 6613 24903 6647
rect 26525 6613 26559 6647
rect 1593 6409 1627 6443
rect 5917 6409 5951 6443
rect 6193 6409 6227 6443
rect 7757 6409 7791 6443
rect 9137 6409 9171 6443
rect 11989 6409 12023 6443
rect 12449 6409 12483 6443
rect 14013 6409 14047 6443
rect 17693 6409 17727 6443
rect 19533 6409 19567 6443
rect 22385 6409 22419 6443
rect 25145 6409 25179 6443
rect 6622 6341 6656 6375
rect 19253 6341 19287 6375
rect 22017 6341 22051 6375
rect 23940 6341 23974 6375
rect 25605 6341 25639 6375
rect 1409 6273 1443 6307
rect 5733 6273 5767 6307
rect 6009 6273 6043 6307
rect 8401 6273 8435 6307
rect 8585 6273 8619 6307
rect 8769 6273 8803 6307
rect 8861 6273 8895 6307
rect 8953 6273 8987 6307
rect 11897 6273 11931 6307
rect 12357 6273 12391 6307
rect 12817 6273 12851 6307
rect 13829 6273 13863 6307
rect 17601 6273 17635 6307
rect 18061 6273 18095 6307
rect 18981 6273 19015 6307
rect 19165 6273 19199 6307
rect 19395 6273 19429 6307
rect 21833 6273 21867 6307
rect 22109 6273 22143 6307
rect 22201 6273 22235 6307
rect 25513 6273 25547 6307
rect 25973 6273 26007 6307
rect 6377 6205 6411 6239
rect 12541 6205 12575 6239
rect 13369 6205 13403 6239
rect 17877 6205 17911 6239
rect 18613 6205 18647 6239
rect 21557 6205 21591 6239
rect 23673 6205 23707 6239
rect 25697 6205 25731 6239
rect 26525 6205 26559 6239
rect 25053 6137 25087 6171
rect 7849 6069 7883 6103
rect 11713 6069 11747 6103
rect 17233 6069 17267 6103
rect 21005 6069 21039 6103
rect 6193 5865 6227 5899
rect 12817 5865 12851 5899
rect 18245 5865 18279 5899
rect 23949 5865 23983 5899
rect 25789 5797 25823 5831
rect 6837 5729 6871 5763
rect 11437 5729 11471 5763
rect 14657 5729 14691 5763
rect 16865 5729 16899 5763
rect 18797 5729 18831 5763
rect 18981 5729 19015 5763
rect 20637 5729 20671 5763
rect 20821 5729 20855 5763
rect 21741 5729 21775 5763
rect 21925 5729 21959 5763
rect 24409 5729 24443 5763
rect 6561 5661 6595 5695
rect 15485 5661 15519 5695
rect 19901 5661 19935 5695
rect 20545 5661 20579 5695
rect 24133 5661 24167 5695
rect 6653 5593 6687 5627
rect 11704 5593 11738 5627
rect 14473 5593 14507 5627
rect 14933 5593 14967 5627
rect 17132 5593 17166 5627
rect 18705 5593 18739 5627
rect 19257 5593 19291 5627
rect 24654 5593 24688 5627
rect 14105 5525 14139 5559
rect 14565 5525 14599 5559
rect 18337 5525 18371 5559
rect 20177 5525 20211 5559
rect 21281 5525 21315 5559
rect 21649 5525 21683 5559
rect 8125 5321 8159 5355
rect 8769 5321 8803 5355
rect 14197 5321 14231 5355
rect 17141 5321 17175 5355
rect 18889 5321 18923 5355
rect 19809 5321 19843 5355
rect 21925 5321 21959 5355
rect 20146 5253 20180 5287
rect 8033 5185 8067 5219
rect 8861 5185 8895 5219
rect 9321 5185 9355 5219
rect 13084 5185 13118 5219
rect 17325 5185 17359 5219
rect 17509 5185 17543 5219
rect 17776 5185 17810 5219
rect 19625 5185 19659 5219
rect 19901 5185 19935 5219
rect 21557 5185 21591 5219
rect 22477 5185 22511 5219
rect 8309 5117 8343 5151
rect 8677 5117 8711 5151
rect 9873 5117 9907 5151
rect 12817 5117 12851 5151
rect 21281 5049 21315 5083
rect 7665 4981 7699 5015
rect 9229 4981 9263 5015
rect 21373 4981 21407 5015
rect 8953 4777 8987 4811
rect 13185 4777 13219 4811
rect 17877 4777 17911 4811
rect 22109 4777 22143 4811
rect 8769 4709 8803 4743
rect 7389 4641 7423 4675
rect 15577 4641 15611 4675
rect 20729 4641 20763 4675
rect 7113 4573 7147 4607
rect 9505 4573 9539 4607
rect 9873 4573 9907 4607
rect 11069 4573 11103 4607
rect 13369 4573 13403 4607
rect 15301 4573 15335 4607
rect 18061 4573 18095 4607
rect 20996 4573 21030 4607
rect 7656 4505 7690 4539
rect 7297 4437 7331 4471
rect 9689 4437 9723 4471
rect 10517 4437 10551 4471
rect 17049 4437 17083 4471
rect 8493 4233 8527 4267
rect 10057 4233 10091 4267
rect 15025 4233 15059 4267
rect 7380 4165 7414 4199
rect 10885 4165 10919 4199
rect 11529 4165 11563 4199
rect 15853 4165 15887 4199
rect 7113 4097 7147 4131
rect 10149 4097 10183 4131
rect 10977 4097 11011 4131
rect 14933 4097 14967 4131
rect 10241 4029 10275 4063
rect 11069 4029 11103 4063
rect 12081 4029 12115 4063
rect 14749 4029 14783 4063
rect 15945 4029 15979 4063
rect 16037 4029 16071 4063
rect 9689 3893 9723 3927
rect 10517 3893 10551 3927
rect 15393 3893 15427 3927
rect 15485 3893 15519 3927
rect 17417 3689 17451 3723
rect 15301 3621 15335 3655
rect 12173 3553 12207 3587
rect 14565 3553 14599 3587
rect 14657 3553 14691 3587
rect 15669 3553 15703 3587
rect 9689 3485 9723 3519
rect 9965 3485 9999 3519
rect 10057 3485 10091 3519
rect 10333 3485 10367 3519
rect 15117 3485 15151 3519
rect 15393 3485 15427 3519
rect 10609 3417 10643 3451
rect 12449 3417 12483 3451
rect 14473 3417 14507 3451
rect 15945 3417 15979 3451
rect 9505 3349 9539 3383
rect 9873 3349 9907 3383
rect 10241 3349 10275 3383
rect 12081 3349 12115 3383
rect 13921 3349 13955 3383
rect 14105 3349 14139 3383
rect 15577 3349 15611 3383
rect 10793 3145 10827 3179
rect 11621 3145 11655 3179
rect 13093 3145 13127 3179
rect 13737 3145 13771 3179
rect 16313 3145 16347 3179
rect 16773 3145 16807 3179
rect 9321 3077 9355 3111
rect 9045 3009 9079 3043
rect 11713 3009 11747 3043
rect 13277 3009 13311 3043
rect 13829 3009 13863 3043
rect 16221 3009 16255 3043
rect 16681 3009 16715 3043
rect 29285 2601 29319 2635
rect 1777 2397 1811 2431
rect 11897 2397 11931 2431
rect 17601 2397 17635 2431
rect 23397 2397 23431 2431
rect 29101 2397 29135 2431
rect 31217 2397 31251 2431
rect 1409 2329 1443 2363
rect 6101 2329 6135 2363
rect 5825 2261 5859 2295
rect 11621 2261 11655 2295
rect 17693 2261 17727 2295
rect 23489 2261 23523 2295
rect 31401 2261 31435 2295
<< metal1 >>
rect 1104 32666 31832 32688
rect 1104 32614 4922 32666
rect 4974 32614 4986 32666
rect 5038 32614 5050 32666
rect 5102 32614 5114 32666
rect 5166 32614 5178 32666
rect 5230 32614 5242 32666
rect 5294 32614 10922 32666
rect 10974 32614 10986 32666
rect 11038 32614 11050 32666
rect 11102 32614 11114 32666
rect 11166 32614 11178 32666
rect 11230 32614 11242 32666
rect 11294 32614 16922 32666
rect 16974 32614 16986 32666
rect 17038 32614 17050 32666
rect 17102 32614 17114 32666
rect 17166 32614 17178 32666
rect 17230 32614 17242 32666
rect 17294 32614 22922 32666
rect 22974 32614 22986 32666
rect 23038 32614 23050 32666
rect 23102 32614 23114 32666
rect 23166 32614 23178 32666
rect 23230 32614 23242 32666
rect 23294 32614 28922 32666
rect 28974 32614 28986 32666
rect 29038 32614 29050 32666
rect 29102 32614 29114 32666
rect 29166 32614 29178 32666
rect 29230 32614 29242 32666
rect 29294 32614 31832 32666
rect 1104 32592 31832 32614
rect 1302 32512 1308 32564
rect 1360 32512 1366 32564
rect 18690 32512 18696 32564
rect 18748 32552 18754 32564
rect 19429 32555 19487 32561
rect 19429 32552 19441 32555
rect 18748 32524 19441 32552
rect 18748 32512 18754 32524
rect 19429 32521 19441 32524
rect 19475 32521 19487 32555
rect 19429 32515 19487 32521
rect 24486 32512 24492 32564
rect 24544 32552 24550 32564
rect 24949 32555 25007 32561
rect 24949 32552 24961 32555
rect 24544 32524 24961 32552
rect 24544 32512 24550 32524
rect 24949 32521 24961 32524
rect 24995 32521 25007 32555
rect 24949 32515 25007 32521
rect 1320 32416 1348 32512
rect 1397 32419 1455 32425
rect 1397 32416 1409 32419
rect 1320 32388 1409 32416
rect 1397 32385 1409 32388
rect 1443 32385 1455 32419
rect 1397 32379 1455 32385
rect 7098 32376 7104 32428
rect 7156 32416 7162 32428
rect 7193 32419 7251 32425
rect 7193 32416 7205 32419
rect 7156 32388 7205 32416
rect 7156 32376 7162 32388
rect 7193 32385 7205 32388
rect 7239 32385 7251 32419
rect 7193 32379 7251 32385
rect 12894 32376 12900 32428
rect 12952 32416 12958 32428
rect 12989 32419 13047 32425
rect 12989 32416 13001 32419
rect 12952 32388 13001 32416
rect 12952 32376 12958 32388
rect 12989 32385 13001 32388
rect 13035 32385 13047 32419
rect 12989 32379 13047 32385
rect 19334 32376 19340 32428
rect 19392 32376 19398 32428
rect 24670 32376 24676 32428
rect 24728 32376 24734 32428
rect 30282 32376 30288 32428
rect 30340 32416 30346 32428
rect 30377 32419 30435 32425
rect 30377 32416 30389 32419
rect 30340 32388 30389 32416
rect 30340 32376 30346 32388
rect 30377 32385 30389 32388
rect 30423 32385 30435 32419
rect 30377 32379 30435 32385
rect 1581 32283 1639 32289
rect 1581 32249 1593 32283
rect 1627 32280 1639 32283
rect 12434 32280 12440 32292
rect 1627 32252 12440 32280
rect 1627 32249 1639 32252
rect 1581 32243 1639 32249
rect 12434 32240 12440 32252
rect 12492 32240 12498 32292
rect 7374 32172 7380 32224
rect 7432 32172 7438 32224
rect 13170 32172 13176 32224
rect 13228 32172 13234 32224
rect 30558 32172 30564 32224
rect 30616 32172 30622 32224
rect 1104 32122 31832 32144
rect 1104 32070 4182 32122
rect 4234 32070 4246 32122
rect 4298 32070 4310 32122
rect 4362 32070 4374 32122
rect 4426 32070 4438 32122
rect 4490 32070 4502 32122
rect 4554 32070 10182 32122
rect 10234 32070 10246 32122
rect 10298 32070 10310 32122
rect 10362 32070 10374 32122
rect 10426 32070 10438 32122
rect 10490 32070 10502 32122
rect 10554 32070 16182 32122
rect 16234 32070 16246 32122
rect 16298 32070 16310 32122
rect 16362 32070 16374 32122
rect 16426 32070 16438 32122
rect 16490 32070 16502 32122
rect 16554 32070 22182 32122
rect 22234 32070 22246 32122
rect 22298 32070 22310 32122
rect 22362 32070 22374 32122
rect 22426 32070 22438 32122
rect 22490 32070 22502 32122
rect 22554 32070 28182 32122
rect 28234 32070 28246 32122
rect 28298 32070 28310 32122
rect 28362 32070 28374 32122
rect 28426 32070 28438 32122
rect 28490 32070 28502 32122
rect 28554 32070 31832 32122
rect 1104 32048 31832 32070
rect 19889 31807 19947 31813
rect 19889 31773 19901 31807
rect 19935 31804 19947 31807
rect 20162 31804 20168 31816
rect 19935 31776 20168 31804
rect 19935 31773 19947 31776
rect 19889 31767 19947 31773
rect 20162 31764 20168 31776
rect 20220 31764 20226 31816
rect 13538 31696 13544 31748
rect 13596 31736 13602 31748
rect 13596 31708 19380 31736
rect 13596 31696 13602 31708
rect 19352 31680 19380 31708
rect 18230 31628 18236 31680
rect 18288 31668 18294 31680
rect 19245 31671 19303 31677
rect 19245 31668 19257 31671
rect 18288 31640 19257 31668
rect 18288 31628 18294 31640
rect 19245 31637 19257 31640
rect 19291 31637 19303 31671
rect 19245 31631 19303 31637
rect 19334 31628 19340 31680
rect 19392 31628 19398 31680
rect 1104 31578 31832 31600
rect 1104 31526 4922 31578
rect 4974 31526 4986 31578
rect 5038 31526 5050 31578
rect 5102 31526 5114 31578
rect 5166 31526 5178 31578
rect 5230 31526 5242 31578
rect 5294 31526 10922 31578
rect 10974 31526 10986 31578
rect 11038 31526 11050 31578
rect 11102 31526 11114 31578
rect 11166 31526 11178 31578
rect 11230 31526 11242 31578
rect 11294 31526 16922 31578
rect 16974 31526 16986 31578
rect 17038 31526 17050 31578
rect 17102 31526 17114 31578
rect 17166 31526 17178 31578
rect 17230 31526 17242 31578
rect 17294 31526 22922 31578
rect 22974 31526 22986 31578
rect 23038 31526 23050 31578
rect 23102 31526 23114 31578
rect 23166 31526 23178 31578
rect 23230 31526 23242 31578
rect 23294 31526 28922 31578
rect 28974 31526 28986 31578
rect 29038 31526 29050 31578
rect 29102 31526 29114 31578
rect 29166 31526 29178 31578
rect 29230 31526 29242 31578
rect 29294 31526 31832 31578
rect 1104 31504 31832 31526
rect 13538 31424 13544 31476
rect 13596 31424 13602 31476
rect 15565 31467 15623 31473
rect 13648 31436 14412 31464
rect 11977 31331 12035 31337
rect 11977 31297 11989 31331
rect 12023 31328 12035 31331
rect 12345 31331 12403 31337
rect 12345 31328 12357 31331
rect 12023 31300 12357 31328
rect 12023 31297 12035 31300
rect 11977 31291 12035 31297
rect 12345 31297 12357 31300
rect 12391 31297 12403 31331
rect 12345 31291 12403 31297
rect 13265 31331 13323 31337
rect 13265 31297 13277 31331
rect 13311 31328 13323 31331
rect 13648 31328 13676 31436
rect 14384 31408 14412 31436
rect 15565 31433 15577 31467
rect 15611 31464 15623 31467
rect 24670 31464 24676 31476
rect 15611 31436 24676 31464
rect 15611 31433 15623 31436
rect 15565 31427 15623 31433
rect 24670 31424 24676 31436
rect 24728 31424 24734 31476
rect 13998 31396 14004 31408
rect 13740 31368 14004 31396
rect 13740 31337 13768 31368
rect 13998 31356 14004 31368
rect 14056 31356 14062 31408
rect 14366 31356 14372 31408
rect 14424 31356 14430 31408
rect 14826 31356 14832 31408
rect 14884 31356 14890 31408
rect 17681 31399 17739 31405
rect 16776 31368 17632 31396
rect 16776 31340 16804 31368
rect 13311 31300 13676 31328
rect 13725 31331 13783 31337
rect 13311 31297 13323 31300
rect 13265 31291 13323 31297
rect 13725 31297 13737 31331
rect 13771 31297 13783 31331
rect 13725 31291 13783 31297
rect 16758 31288 16764 31340
rect 16816 31288 16822 31340
rect 17052 31337 17080 31368
rect 16945 31331 17003 31337
rect 16945 31297 16957 31331
rect 16991 31297 17003 31331
rect 16945 31291 17003 31297
rect 17037 31331 17095 31337
rect 17037 31297 17049 31331
rect 17083 31297 17095 31331
rect 17037 31291 17095 31297
rect 17129 31331 17187 31337
rect 17129 31297 17141 31331
rect 17175 31328 17187 31331
rect 17218 31328 17224 31340
rect 17175 31300 17224 31328
rect 17175 31297 17187 31300
rect 17129 31291 17187 31297
rect 10778 31220 10784 31272
rect 10836 31220 10842 31272
rect 12069 31263 12127 31269
rect 12069 31229 12081 31263
rect 12115 31260 12127 31263
rect 12802 31260 12808 31272
rect 12115 31232 12808 31260
rect 12115 31229 12127 31232
rect 12069 31223 12127 31229
rect 12802 31220 12808 31232
rect 12860 31220 12866 31272
rect 12894 31220 12900 31272
rect 12952 31220 12958 31272
rect 13817 31263 13875 31269
rect 13817 31229 13829 31263
rect 13863 31229 13875 31263
rect 13817 31223 13875 31229
rect 10796 31192 10824 31220
rect 13832 31192 13860 31223
rect 14090 31220 14096 31272
rect 14148 31220 14154 31272
rect 10796 31164 13860 31192
rect 16960 31192 16988 31291
rect 17218 31288 17224 31300
rect 17276 31288 17282 31340
rect 17420 31337 17448 31368
rect 17313 31331 17371 31337
rect 17313 31297 17325 31331
rect 17359 31297 17371 31331
rect 17313 31291 17371 31297
rect 17405 31331 17463 31337
rect 17405 31297 17417 31331
rect 17451 31297 17463 31331
rect 17405 31291 17463 31297
rect 17328 31260 17356 31291
rect 17494 31288 17500 31340
rect 17552 31288 17558 31340
rect 17604 31328 17632 31368
rect 17681 31365 17693 31399
rect 17727 31396 17739 31399
rect 18230 31396 18236 31408
rect 17727 31368 18236 31396
rect 17727 31365 17739 31368
rect 17681 31359 17739 31365
rect 18230 31356 18236 31368
rect 18288 31356 18294 31408
rect 18693 31399 18751 31405
rect 18693 31396 18705 31399
rect 18340 31368 18705 31396
rect 17773 31331 17831 31337
rect 17773 31328 17785 31331
rect 17604 31300 17785 31328
rect 17773 31297 17785 31300
rect 17819 31297 17831 31331
rect 17773 31291 17831 31297
rect 17862 31288 17868 31340
rect 17920 31288 17926 31340
rect 18049 31331 18107 31337
rect 18049 31328 18061 31331
rect 17972 31300 18061 31328
rect 17586 31260 17592 31272
rect 17328 31232 17592 31260
rect 17586 31220 17592 31232
rect 17644 31220 17650 31272
rect 17972 31260 18000 31300
rect 18049 31297 18061 31300
rect 18095 31297 18107 31331
rect 18049 31291 18107 31297
rect 18340 31260 18368 31368
rect 18693 31365 18705 31368
rect 18739 31365 18751 31399
rect 18693 31359 18751 31365
rect 19426 31356 19432 31408
rect 19484 31356 19490 31408
rect 17696 31232 18000 31260
rect 18064 31232 18368 31260
rect 18417 31263 18475 31269
rect 17696 31201 17724 31232
rect 18064 31201 18092 31232
rect 18417 31229 18429 31263
rect 18463 31260 18475 31263
rect 18782 31260 18788 31272
rect 18463 31232 18788 31260
rect 18463 31229 18475 31232
rect 18417 31223 18475 31229
rect 18782 31220 18788 31232
rect 18840 31220 18846 31272
rect 17681 31195 17739 31201
rect 16960 31164 17632 31192
rect 11606 31084 11612 31136
rect 11664 31084 11670 31136
rect 13170 31084 13176 31136
rect 13228 31084 13234 31136
rect 13832 31124 13860 31164
rect 15470 31124 15476 31136
rect 13832 31096 15476 31124
rect 15470 31084 15476 31096
rect 15528 31084 15534 31136
rect 16850 31084 16856 31136
rect 16908 31084 16914 31136
rect 17310 31084 17316 31136
rect 17368 31084 17374 31136
rect 17604 31124 17632 31164
rect 17681 31161 17693 31195
rect 17727 31161 17739 31195
rect 17681 31155 17739 31161
rect 18049 31195 18107 31201
rect 18049 31161 18061 31195
rect 18095 31161 18107 31195
rect 18049 31155 18107 31161
rect 20162 31152 20168 31204
rect 20220 31152 20226 31204
rect 17770 31124 17776 31136
rect 17604 31096 17776 31124
rect 17770 31084 17776 31096
rect 17828 31124 17834 31136
rect 18506 31124 18512 31136
rect 17828 31096 18512 31124
rect 17828 31084 17834 31096
rect 18506 31084 18512 31096
rect 18564 31084 18570 31136
rect 1104 31034 31832 31056
rect 1104 30982 4182 31034
rect 4234 30982 4246 31034
rect 4298 30982 4310 31034
rect 4362 30982 4374 31034
rect 4426 30982 4438 31034
rect 4490 30982 4502 31034
rect 4554 30982 10182 31034
rect 10234 30982 10246 31034
rect 10298 30982 10310 31034
rect 10362 30982 10374 31034
rect 10426 30982 10438 31034
rect 10490 30982 10502 31034
rect 10554 30982 16182 31034
rect 16234 30982 16246 31034
rect 16298 30982 16310 31034
rect 16362 30982 16374 31034
rect 16426 30982 16438 31034
rect 16490 30982 16502 31034
rect 16554 30982 22182 31034
rect 22234 30982 22246 31034
rect 22298 30982 22310 31034
rect 22362 30982 22374 31034
rect 22426 30982 22438 31034
rect 22490 30982 22502 31034
rect 22554 30982 28182 31034
rect 28234 30982 28246 31034
rect 28298 30982 28310 31034
rect 28362 30982 28374 31034
rect 28426 30982 28438 31034
rect 28490 30982 28502 31034
rect 28554 30982 31832 31034
rect 1104 30960 31832 30982
rect 13170 30920 13176 30932
rect 12406 30892 13176 30920
rect 11057 30787 11115 30793
rect 11057 30753 11069 30787
rect 11103 30784 11115 30787
rect 11606 30784 11612 30796
rect 11103 30756 11612 30784
rect 11103 30753 11115 30756
rect 11057 30747 11115 30753
rect 11606 30744 11612 30756
rect 11664 30744 11670 30796
rect 12406 30784 12434 30892
rect 13170 30880 13176 30892
rect 13228 30880 13234 30932
rect 13538 30880 13544 30932
rect 13596 30880 13602 30932
rect 13725 30923 13783 30929
rect 13725 30889 13737 30923
rect 13771 30920 13783 30923
rect 14090 30920 14096 30932
rect 13771 30892 14096 30920
rect 13771 30889 13783 30892
rect 13725 30883 13783 30889
rect 14090 30880 14096 30892
rect 14148 30880 14154 30932
rect 14826 30880 14832 30932
rect 14884 30880 14890 30932
rect 17310 30880 17316 30932
rect 17368 30880 17374 30932
rect 17586 30880 17592 30932
rect 17644 30920 17650 30932
rect 18417 30923 18475 30929
rect 18417 30920 18429 30923
rect 17644 30892 18429 30920
rect 17644 30880 17650 30892
rect 18417 30889 18429 30892
rect 18463 30889 18475 30923
rect 21005 30923 21063 30929
rect 21005 30920 21017 30923
rect 18417 30883 18475 30889
rect 19628 30892 21017 30920
rect 12529 30855 12587 30861
rect 12529 30821 12541 30855
rect 12575 30852 12587 30855
rect 12894 30852 12900 30864
rect 12575 30824 12900 30852
rect 12575 30821 12587 30824
rect 12529 30815 12587 30821
rect 12894 30812 12900 30824
rect 12952 30812 12958 30864
rect 12176 30756 12434 30784
rect 934 30676 940 30728
rect 992 30716 998 30728
rect 1397 30719 1455 30725
rect 1397 30716 1409 30719
rect 992 30688 1409 30716
rect 992 30676 998 30688
rect 1397 30685 1409 30688
rect 1443 30685 1455 30719
rect 1397 30679 1455 30685
rect 10778 30676 10784 30728
rect 10836 30676 10842 30728
rect 12176 30702 12204 30756
rect 12434 30676 12440 30728
rect 12492 30716 12498 30728
rect 12986 30716 12992 30728
rect 12492 30688 12992 30716
rect 12492 30676 12498 30688
rect 12986 30676 12992 30688
rect 13044 30716 13050 30728
rect 13556 30725 13584 30880
rect 15470 30744 15476 30796
rect 15528 30744 15534 30796
rect 17328 30784 17356 30880
rect 18325 30855 18383 30861
rect 18325 30821 18337 30855
rect 18371 30852 18383 30855
rect 19628 30852 19656 30892
rect 21005 30889 21017 30892
rect 21051 30889 21063 30923
rect 21005 30883 21063 30889
rect 18371 30824 19656 30852
rect 18371 30821 18383 30824
rect 18325 30815 18383 30821
rect 21269 30787 21327 30793
rect 21269 30784 21281 30787
rect 17328 30756 18368 30784
rect 13173 30719 13231 30725
rect 13173 30716 13185 30719
rect 13044 30688 13185 30716
rect 13044 30676 13050 30688
rect 13173 30685 13185 30688
rect 13219 30685 13231 30719
rect 13173 30679 13231 30685
rect 13541 30719 13599 30725
rect 13541 30685 13553 30719
rect 13587 30685 13599 30719
rect 13541 30679 13599 30685
rect 14277 30719 14335 30725
rect 14277 30685 14289 30719
rect 14323 30685 14335 30719
rect 14737 30719 14795 30725
rect 14737 30716 14749 30719
rect 14277 30679 14335 30685
rect 14384 30688 14749 30716
rect 13357 30651 13415 30657
rect 13357 30617 13369 30651
rect 13403 30617 13415 30651
rect 13357 30611 13415 30617
rect 1578 30540 1584 30592
rect 1636 30540 1642 30592
rect 13372 30580 13400 30611
rect 13446 30608 13452 30660
rect 13504 30608 13510 30660
rect 14090 30608 14096 30660
rect 14148 30608 14154 30660
rect 14108 30580 14136 30608
rect 14292 30592 14320 30679
rect 14384 30592 14412 30688
rect 14737 30685 14749 30688
rect 14783 30716 14795 30719
rect 15010 30716 15016 30728
rect 14783 30688 15016 30716
rect 14783 30685 14795 30688
rect 14737 30679 14795 30685
rect 15010 30676 15016 30688
rect 15068 30676 15074 30728
rect 16850 30676 16856 30728
rect 16908 30676 16914 30728
rect 17957 30719 18015 30725
rect 17957 30716 17969 30719
rect 17236 30688 17969 30716
rect 15746 30608 15752 30660
rect 15804 30608 15810 30660
rect 13372 30552 14136 30580
rect 14182 30540 14188 30592
rect 14240 30540 14246 30592
rect 14274 30540 14280 30592
rect 14332 30540 14338 30592
rect 14366 30540 14372 30592
rect 14424 30540 14430 30592
rect 16574 30540 16580 30592
rect 16632 30580 16638 30592
rect 17236 30589 17264 30688
rect 17957 30685 17969 30688
rect 18003 30685 18015 30719
rect 17957 30679 18015 30685
rect 18138 30676 18144 30728
rect 18196 30676 18202 30728
rect 18340 30725 18368 30756
rect 18800 30756 21281 30784
rect 18800 30728 18828 30756
rect 21269 30753 21281 30756
rect 21315 30753 21327 30787
rect 21269 30747 21327 30753
rect 18325 30719 18383 30725
rect 18325 30685 18337 30719
rect 18371 30685 18383 30719
rect 18325 30679 18383 30685
rect 18782 30676 18788 30728
rect 18840 30676 18846 30728
rect 19061 30719 19119 30725
rect 19061 30685 19073 30719
rect 19107 30716 19119 30719
rect 19245 30719 19303 30725
rect 19245 30716 19257 30719
rect 19107 30688 19257 30716
rect 19107 30685 19119 30688
rect 19061 30679 19119 30685
rect 19245 30685 19257 30688
rect 19291 30716 19303 30719
rect 19334 30716 19340 30728
rect 19291 30688 19340 30716
rect 19291 30685 19303 30688
rect 19245 30679 19303 30685
rect 17310 30608 17316 30660
rect 17368 30648 17374 30660
rect 17862 30648 17868 30660
rect 17368 30620 17868 30648
rect 17368 30608 17374 30620
rect 17862 30608 17868 30620
rect 17920 30608 17926 30660
rect 17221 30583 17279 30589
rect 17221 30580 17233 30583
rect 16632 30552 17233 30580
rect 16632 30540 16638 30552
rect 17221 30549 17233 30552
rect 17267 30549 17279 30583
rect 17221 30543 17279 30549
rect 17402 30540 17408 30592
rect 17460 30540 17466 30592
rect 17586 30540 17592 30592
rect 17644 30580 17650 30592
rect 19076 30580 19104 30679
rect 19334 30676 19340 30688
rect 19392 30676 19398 30728
rect 19518 30608 19524 30660
rect 19576 30648 19582 30660
rect 19576 30620 19826 30648
rect 19576 30608 19582 30620
rect 17644 30552 19104 30580
rect 17644 30540 17650 30552
rect 1104 30490 31832 30512
rect 1104 30438 4922 30490
rect 4974 30438 4986 30490
rect 5038 30438 5050 30490
rect 5102 30438 5114 30490
rect 5166 30438 5178 30490
rect 5230 30438 5242 30490
rect 5294 30438 10922 30490
rect 10974 30438 10986 30490
rect 11038 30438 11050 30490
rect 11102 30438 11114 30490
rect 11166 30438 11178 30490
rect 11230 30438 11242 30490
rect 11294 30438 16922 30490
rect 16974 30438 16986 30490
rect 17038 30438 17050 30490
rect 17102 30438 17114 30490
rect 17166 30438 17178 30490
rect 17230 30438 17242 30490
rect 17294 30438 22922 30490
rect 22974 30438 22986 30490
rect 23038 30438 23050 30490
rect 23102 30438 23114 30490
rect 23166 30438 23178 30490
rect 23230 30438 23242 30490
rect 23294 30438 28922 30490
rect 28974 30438 28986 30490
rect 29038 30438 29050 30490
rect 29102 30438 29114 30490
rect 29166 30438 29178 30490
rect 29230 30438 29242 30490
rect 29294 30438 31832 30490
rect 1104 30416 31832 30438
rect 12802 30336 12808 30388
rect 12860 30336 12866 30388
rect 15657 30379 15715 30385
rect 15657 30345 15669 30379
rect 15703 30376 15715 30379
rect 15746 30376 15752 30388
rect 15703 30348 15752 30376
rect 15703 30345 15715 30348
rect 15657 30339 15715 30345
rect 15746 30336 15752 30348
rect 15804 30336 15810 30388
rect 15841 30379 15899 30385
rect 15841 30345 15853 30379
rect 15887 30345 15899 30379
rect 15841 30339 15899 30345
rect 18248 30348 19104 30376
rect 12820 30308 12848 30336
rect 14737 30311 14795 30317
rect 14737 30308 14749 30311
rect 12820 30280 14749 30308
rect 14737 30277 14749 30280
rect 14783 30308 14795 30311
rect 15856 30308 15884 30339
rect 16666 30308 16672 30320
rect 14783 30280 15884 30308
rect 16132 30280 16672 30308
rect 14783 30277 14795 30280
rect 14737 30271 14795 30277
rect 11882 30200 11888 30252
rect 11940 30200 11946 30252
rect 12621 30243 12679 30249
rect 12621 30209 12633 30243
rect 12667 30240 12679 30243
rect 12894 30240 12900 30252
rect 12667 30212 12900 30240
rect 12667 30209 12679 30212
rect 12621 30203 12679 30209
rect 12894 30200 12900 30212
rect 12952 30200 12958 30252
rect 13906 30200 13912 30252
rect 13964 30200 13970 30252
rect 14918 30200 14924 30252
rect 14976 30200 14982 30252
rect 15010 30200 15016 30252
rect 15068 30240 15074 30252
rect 15068 30212 15240 30240
rect 15068 30200 15074 30212
rect 14642 30132 14648 30184
rect 14700 30172 14706 30184
rect 15105 30175 15163 30181
rect 15105 30172 15117 30175
rect 14700 30144 15117 30172
rect 14700 30132 14706 30144
rect 15105 30141 15117 30144
rect 15151 30141 15163 30175
rect 15105 30135 15163 30141
rect 13541 30039 13599 30045
rect 13541 30005 13553 30039
rect 13587 30036 13599 30039
rect 13630 30036 13636 30048
rect 13587 30008 13636 30036
rect 13587 30005 13599 30008
rect 13541 29999 13599 30005
rect 13630 29996 13636 30008
rect 13688 29996 13694 30048
rect 14001 30039 14059 30045
rect 14001 30005 14013 30039
rect 14047 30036 14059 30039
rect 14090 30036 14096 30048
rect 14047 30008 14096 30036
rect 14047 30005 14059 30008
rect 14001 29999 14059 30005
rect 14090 29996 14096 30008
rect 14148 29996 14154 30048
rect 15120 30036 15148 30135
rect 15212 30104 15240 30212
rect 15746 30200 15752 30252
rect 15804 30249 15810 30252
rect 15804 30243 15840 30249
rect 15828 30209 15840 30243
rect 15804 30203 15840 30209
rect 15804 30200 15810 30203
rect 16132 30172 16160 30280
rect 16666 30268 16672 30280
rect 16724 30308 16730 30320
rect 16724 30280 18184 30308
rect 16724 30268 16730 30280
rect 18156 30252 18184 30280
rect 16209 30243 16267 30249
rect 16209 30209 16221 30243
rect 16255 30240 16267 30243
rect 17402 30240 17408 30252
rect 16255 30212 17408 30240
rect 16255 30209 16267 30212
rect 16209 30203 16267 30209
rect 17402 30200 17408 30212
rect 17460 30200 17466 30252
rect 17494 30200 17500 30252
rect 17552 30200 17558 30252
rect 17589 30243 17647 30249
rect 17589 30209 17601 30243
rect 17635 30240 17647 30243
rect 17770 30240 17776 30252
rect 17635 30212 17776 30240
rect 17635 30209 17647 30212
rect 17589 30203 17647 30209
rect 17770 30200 17776 30212
rect 17828 30200 17834 30252
rect 17865 30243 17923 30249
rect 17865 30209 17877 30243
rect 17911 30209 17923 30243
rect 17865 30203 17923 30209
rect 16301 30175 16359 30181
rect 16301 30172 16313 30175
rect 16132 30144 16313 30172
rect 16301 30141 16313 30144
rect 16347 30141 16359 30175
rect 16301 30135 16359 30141
rect 16761 30175 16819 30181
rect 16761 30141 16773 30175
rect 16807 30141 16819 30175
rect 17512 30172 17540 30200
rect 17880 30172 17908 30203
rect 18138 30200 18144 30252
rect 18196 30200 18202 30252
rect 18248 30181 18276 30348
rect 19076 30317 19104 30348
rect 19061 30311 19119 30317
rect 19061 30277 19073 30311
rect 19107 30277 19119 30311
rect 19061 30271 19119 30277
rect 19702 30268 19708 30320
rect 19760 30268 19766 30320
rect 18506 30200 18512 30252
rect 18564 30200 18570 30252
rect 17512 30144 17908 30172
rect 17957 30175 18015 30181
rect 16761 30135 16819 30141
rect 17957 30141 17969 30175
rect 18003 30141 18015 30175
rect 17957 30135 18015 30141
rect 18233 30175 18291 30181
rect 18233 30141 18245 30175
rect 18279 30141 18291 30175
rect 18782 30172 18788 30184
rect 18233 30135 18291 30141
rect 18524 30144 18788 30172
rect 16776 30104 16804 30135
rect 17972 30104 18000 30135
rect 15212 30076 16804 30104
rect 17880 30076 18000 30104
rect 16758 30036 16764 30048
rect 15120 30008 16764 30036
rect 16758 29996 16764 30008
rect 16816 29996 16822 30048
rect 16850 29996 16856 30048
rect 16908 30036 16914 30048
rect 17880 30036 17908 30076
rect 16908 30008 17908 30036
rect 16908 29996 16914 30008
rect 17954 29996 17960 30048
rect 18012 30036 18018 30048
rect 18524 30036 18552 30144
rect 18782 30132 18788 30144
rect 18840 30132 18846 30184
rect 19518 30172 19524 30184
rect 18892 30144 19524 30172
rect 18012 30008 18552 30036
rect 18601 30039 18659 30045
rect 18012 29996 18018 30008
rect 18601 30005 18613 30039
rect 18647 30036 18659 30039
rect 18892 30036 18920 30144
rect 19518 30132 19524 30144
rect 19576 30132 19582 30184
rect 18647 30008 18920 30036
rect 18647 30005 18659 30008
rect 18601 29999 18659 30005
rect 20438 29996 20444 30048
rect 20496 30036 20502 30048
rect 20533 30039 20591 30045
rect 20533 30036 20545 30039
rect 20496 30008 20545 30036
rect 20496 29996 20502 30008
rect 20533 30005 20545 30008
rect 20579 30005 20591 30039
rect 20533 29999 20591 30005
rect 1104 29946 31832 29968
rect 1104 29894 4182 29946
rect 4234 29894 4246 29946
rect 4298 29894 4310 29946
rect 4362 29894 4374 29946
rect 4426 29894 4438 29946
rect 4490 29894 4502 29946
rect 4554 29894 10182 29946
rect 10234 29894 10246 29946
rect 10298 29894 10310 29946
rect 10362 29894 10374 29946
rect 10426 29894 10438 29946
rect 10490 29894 10502 29946
rect 10554 29894 16182 29946
rect 16234 29894 16246 29946
rect 16298 29894 16310 29946
rect 16362 29894 16374 29946
rect 16426 29894 16438 29946
rect 16490 29894 16502 29946
rect 16554 29894 22182 29946
rect 22234 29894 22246 29946
rect 22298 29894 22310 29946
rect 22362 29894 22374 29946
rect 22426 29894 22438 29946
rect 22490 29894 22502 29946
rect 22554 29894 28182 29946
rect 28234 29894 28246 29946
rect 28298 29894 28310 29946
rect 28362 29894 28374 29946
rect 28426 29894 28438 29946
rect 28490 29894 28502 29946
rect 28554 29894 31832 29946
rect 1104 29872 31832 29894
rect 13906 29792 13912 29844
rect 13964 29792 13970 29844
rect 13998 29792 14004 29844
rect 14056 29832 14062 29844
rect 14093 29835 14151 29841
rect 14093 29832 14105 29835
rect 14056 29804 14105 29832
rect 14056 29792 14062 29804
rect 14093 29801 14105 29804
rect 14139 29801 14151 29835
rect 14093 29795 14151 29801
rect 14918 29792 14924 29844
rect 14976 29832 14982 29844
rect 16209 29835 16267 29841
rect 16209 29832 16221 29835
rect 14976 29804 16221 29832
rect 14976 29792 14982 29804
rect 16209 29801 16221 29804
rect 16255 29801 16267 29835
rect 16209 29795 16267 29801
rect 16666 29792 16672 29844
rect 16724 29792 16730 29844
rect 16758 29792 16764 29844
rect 16816 29832 16822 29844
rect 16853 29835 16911 29841
rect 16853 29832 16865 29835
rect 16816 29804 16865 29832
rect 16816 29792 16822 29804
rect 16853 29801 16865 29804
rect 16899 29832 16911 29835
rect 17402 29832 17408 29844
rect 16899 29804 17408 29832
rect 16899 29801 16911 29804
rect 16853 29795 16911 29801
rect 17402 29792 17408 29804
rect 17460 29792 17466 29844
rect 17494 29792 17500 29844
rect 17552 29792 17558 29844
rect 19426 29792 19432 29844
rect 19484 29792 19490 29844
rect 19702 29792 19708 29844
rect 19760 29792 19766 29844
rect 15657 29767 15715 29773
rect 13372 29736 14504 29764
rect 12986 29656 12992 29708
rect 13044 29656 13050 29708
rect 13372 29637 13400 29736
rect 13464 29668 13768 29696
rect 13464 29637 13492 29668
rect 13740 29637 13768 29668
rect 13357 29631 13415 29637
rect 13357 29597 13369 29631
rect 13403 29597 13415 29631
rect 13357 29591 13415 29597
rect 13449 29631 13507 29637
rect 13449 29597 13461 29631
rect 13495 29597 13507 29631
rect 13449 29591 13507 29597
rect 13541 29631 13599 29637
rect 13541 29597 13553 29631
rect 13587 29597 13599 29631
rect 13541 29591 13599 29597
rect 13725 29631 13783 29637
rect 13725 29597 13737 29631
rect 13771 29628 13783 29631
rect 14182 29628 14188 29640
rect 13771 29600 14188 29628
rect 13771 29597 13783 29600
rect 13725 29591 13783 29597
rect 13372 29560 13400 29591
rect 13556 29560 13584 29591
rect 14182 29588 14188 29600
rect 14240 29588 14246 29640
rect 14274 29588 14280 29640
rect 14332 29588 14338 29640
rect 14476 29637 14504 29736
rect 15657 29733 15669 29767
rect 15703 29764 15715 29767
rect 16022 29764 16028 29776
rect 15703 29736 16028 29764
rect 15703 29733 15715 29736
rect 15657 29727 15715 29733
rect 16022 29724 16028 29736
rect 16080 29764 16086 29776
rect 17512 29764 17540 29792
rect 16080 29736 17540 29764
rect 16080 29724 16086 29736
rect 15488 29668 16712 29696
rect 15488 29637 15516 29668
rect 14461 29631 14519 29637
rect 14461 29597 14473 29631
rect 14507 29628 14519 29631
rect 15473 29631 15531 29637
rect 14507 29600 15056 29628
rect 14507 29597 14519 29600
rect 14461 29591 14519 29597
rect 14292 29560 14320 29588
rect 13372 29532 13584 29560
rect 13648 29532 14320 29560
rect 13648 29504 13676 29532
rect 15028 29504 15056 29600
rect 15473 29597 15485 29631
rect 15519 29597 15531 29631
rect 15473 29591 15531 29597
rect 16393 29631 16451 29637
rect 16393 29597 16405 29631
rect 16439 29597 16451 29631
rect 16393 29591 16451 29597
rect 16408 29560 16436 29591
rect 16574 29588 16580 29640
rect 16632 29588 16638 29640
rect 16684 29628 16712 29668
rect 17494 29656 17500 29708
rect 17552 29656 17558 29708
rect 18506 29656 18512 29708
rect 18564 29696 18570 29708
rect 18564 29668 19380 29696
rect 18564 29656 18570 29668
rect 17681 29631 17739 29637
rect 17681 29628 17693 29631
rect 16684 29600 17693 29628
rect 17681 29597 17693 29600
rect 17727 29597 17739 29631
rect 17681 29591 17739 29597
rect 17865 29631 17923 29637
rect 17865 29597 17877 29631
rect 17911 29628 17923 29631
rect 18046 29628 18052 29640
rect 17911 29600 18052 29628
rect 17911 29597 17923 29600
rect 17865 29591 17923 29597
rect 17037 29563 17095 29569
rect 17037 29560 17049 29563
rect 16408 29532 17049 29560
rect 17037 29529 17049 29532
rect 17083 29560 17095 29563
rect 17586 29560 17592 29572
rect 17083 29532 17592 29560
rect 17083 29529 17095 29532
rect 17037 29523 17095 29529
rect 17586 29520 17592 29532
rect 17644 29520 17650 29572
rect 17696 29560 17724 29591
rect 18046 29588 18052 29600
rect 18104 29588 18110 29640
rect 19352 29637 19380 29668
rect 19337 29631 19395 29637
rect 19337 29597 19349 29631
rect 19383 29628 19395 29631
rect 19613 29631 19671 29637
rect 19613 29628 19625 29631
rect 19383 29600 19625 29628
rect 19383 29597 19395 29600
rect 19337 29591 19395 29597
rect 19613 29597 19625 29600
rect 19659 29597 19671 29631
rect 19613 29591 19671 29597
rect 20438 29588 20444 29640
rect 20496 29588 20502 29640
rect 20456 29560 20484 29588
rect 17696 29532 20484 29560
rect 13262 29452 13268 29504
rect 13320 29452 13326 29504
rect 13630 29452 13636 29504
rect 13688 29452 13694 29504
rect 15010 29452 15016 29504
rect 15068 29452 15074 29504
rect 15746 29452 15752 29504
rect 15804 29492 15810 29504
rect 16850 29501 16856 29504
rect 16827 29495 16856 29501
rect 16827 29492 16839 29495
rect 15804 29464 16839 29492
rect 15804 29452 15810 29464
rect 16827 29461 16839 29464
rect 16827 29455 16856 29461
rect 16850 29452 16856 29455
rect 16908 29452 16914 29504
rect 17402 29452 17408 29504
rect 17460 29492 17466 29504
rect 17696 29492 17724 29532
rect 17460 29464 17724 29492
rect 17460 29452 17466 29464
rect 1104 29402 31832 29424
rect 1104 29350 4922 29402
rect 4974 29350 4986 29402
rect 5038 29350 5050 29402
rect 5102 29350 5114 29402
rect 5166 29350 5178 29402
rect 5230 29350 5242 29402
rect 5294 29350 10922 29402
rect 10974 29350 10986 29402
rect 11038 29350 11050 29402
rect 11102 29350 11114 29402
rect 11166 29350 11178 29402
rect 11230 29350 11242 29402
rect 11294 29350 16922 29402
rect 16974 29350 16986 29402
rect 17038 29350 17050 29402
rect 17102 29350 17114 29402
rect 17166 29350 17178 29402
rect 17230 29350 17242 29402
rect 17294 29350 22922 29402
rect 22974 29350 22986 29402
rect 23038 29350 23050 29402
rect 23102 29350 23114 29402
rect 23166 29350 23178 29402
rect 23230 29350 23242 29402
rect 23294 29350 28922 29402
rect 28974 29350 28986 29402
rect 29038 29350 29050 29402
rect 29102 29350 29114 29402
rect 29166 29350 29178 29402
rect 29230 29350 29242 29402
rect 29294 29350 31832 29402
rect 1104 29328 31832 29350
rect 13262 29112 13268 29164
rect 13320 29152 13326 29164
rect 13722 29152 13728 29164
rect 13320 29124 13728 29152
rect 13320 29112 13326 29124
rect 13722 29112 13728 29124
rect 13780 29152 13786 29164
rect 14366 29152 14372 29164
rect 13780 29124 14372 29152
rect 13780 29112 13786 29124
rect 14366 29112 14372 29124
rect 14424 29152 14430 29164
rect 14553 29155 14611 29161
rect 14553 29152 14565 29155
rect 14424 29124 14565 29152
rect 14424 29112 14430 29124
rect 14553 29121 14565 29124
rect 14599 29121 14611 29155
rect 14553 29115 14611 29121
rect 15746 29084 15752 29096
rect 14752 29056 15752 29084
rect 14752 29025 14780 29056
rect 15746 29044 15752 29056
rect 15804 29044 15810 29096
rect 14737 29019 14795 29025
rect 14737 28985 14749 29019
rect 14783 28985 14795 29019
rect 14737 28979 14795 28985
rect 1104 28858 31832 28880
rect 1104 28806 4182 28858
rect 4234 28806 4246 28858
rect 4298 28806 4310 28858
rect 4362 28806 4374 28858
rect 4426 28806 4438 28858
rect 4490 28806 4502 28858
rect 4554 28806 10182 28858
rect 10234 28806 10246 28858
rect 10298 28806 10310 28858
rect 10362 28806 10374 28858
rect 10426 28806 10438 28858
rect 10490 28806 10502 28858
rect 10554 28806 16182 28858
rect 16234 28806 16246 28858
rect 16298 28806 16310 28858
rect 16362 28806 16374 28858
rect 16426 28806 16438 28858
rect 16490 28806 16502 28858
rect 16554 28806 22182 28858
rect 22234 28806 22246 28858
rect 22298 28806 22310 28858
rect 22362 28806 22374 28858
rect 22426 28806 22438 28858
rect 22490 28806 22502 28858
rect 22554 28806 28182 28858
rect 28234 28806 28246 28858
rect 28298 28806 28310 28858
rect 28362 28806 28374 28858
rect 28426 28806 28438 28858
rect 28490 28806 28502 28858
rect 28554 28806 31832 28858
rect 1104 28784 31832 28806
rect 11882 28704 11888 28756
rect 11940 28744 11946 28756
rect 12345 28747 12403 28753
rect 12345 28744 12357 28747
rect 11940 28716 12357 28744
rect 11940 28704 11946 28716
rect 12345 28713 12357 28716
rect 12391 28713 12403 28747
rect 12345 28707 12403 28713
rect 8478 28500 8484 28552
rect 8536 28500 8542 28552
rect 8662 28500 8668 28552
rect 8720 28540 8726 28552
rect 8941 28543 8999 28549
rect 8941 28540 8953 28543
rect 8720 28512 8953 28540
rect 8720 28500 8726 28512
rect 8941 28509 8953 28512
rect 8987 28509 8999 28543
rect 8941 28503 8999 28509
rect 10597 28543 10655 28549
rect 10597 28509 10609 28543
rect 10643 28509 10655 28543
rect 10597 28503 10655 28509
rect 9186 28475 9244 28481
rect 9186 28472 9198 28475
rect 8680 28444 9198 28472
rect 8680 28413 8708 28444
rect 9186 28441 9198 28444
rect 9232 28441 9244 28475
rect 10612 28472 10640 28503
rect 14366 28500 14372 28552
rect 14424 28500 14430 28552
rect 14918 28540 14924 28552
rect 14568 28512 14924 28540
rect 10778 28472 10784 28484
rect 10612 28444 10784 28472
rect 9186 28435 9244 28441
rect 10778 28432 10784 28444
rect 10836 28432 10842 28484
rect 10873 28475 10931 28481
rect 10873 28441 10885 28475
rect 10919 28441 10931 28475
rect 12098 28444 12434 28472
rect 10873 28435 10931 28441
rect 8665 28407 8723 28413
rect 8665 28373 8677 28407
rect 8711 28373 8723 28407
rect 8665 28367 8723 28373
rect 10318 28364 10324 28416
rect 10376 28364 10382 28416
rect 10502 28364 10508 28416
rect 10560 28404 10566 28416
rect 10888 28404 10916 28435
rect 10560 28376 10916 28404
rect 12406 28404 12434 28444
rect 13814 28432 13820 28484
rect 13872 28472 13878 28484
rect 14277 28475 14335 28481
rect 13872 28444 14228 28472
rect 13872 28432 13878 28444
rect 13998 28404 14004 28416
rect 12406 28376 14004 28404
rect 10560 28364 10566 28376
rect 13998 28364 14004 28376
rect 14056 28364 14062 28416
rect 14090 28364 14096 28416
rect 14148 28364 14154 28416
rect 14200 28404 14228 28444
rect 14277 28441 14289 28475
rect 14323 28472 14335 28475
rect 14568 28472 14596 28512
rect 14918 28500 14924 28512
rect 14976 28500 14982 28552
rect 14323 28444 14596 28472
rect 14645 28475 14703 28481
rect 14323 28441 14335 28444
rect 14277 28435 14335 28441
rect 14645 28441 14657 28475
rect 14691 28472 14703 28475
rect 14734 28472 14740 28484
rect 14691 28444 14740 28472
rect 14691 28441 14703 28444
rect 14645 28435 14703 28441
rect 14734 28432 14740 28444
rect 14792 28432 14798 28484
rect 14461 28407 14519 28413
rect 14461 28404 14473 28407
rect 14200 28376 14473 28404
rect 14461 28373 14473 28376
rect 14507 28404 14519 28407
rect 14550 28404 14556 28416
rect 14507 28376 14556 28404
rect 14507 28373 14519 28376
rect 14461 28367 14519 28373
rect 14550 28364 14556 28376
rect 14608 28364 14614 28416
rect 1104 28314 31832 28336
rect 1104 28262 4922 28314
rect 4974 28262 4986 28314
rect 5038 28262 5050 28314
rect 5102 28262 5114 28314
rect 5166 28262 5178 28314
rect 5230 28262 5242 28314
rect 5294 28262 10922 28314
rect 10974 28262 10986 28314
rect 11038 28262 11050 28314
rect 11102 28262 11114 28314
rect 11166 28262 11178 28314
rect 11230 28262 11242 28314
rect 11294 28262 16922 28314
rect 16974 28262 16986 28314
rect 17038 28262 17050 28314
rect 17102 28262 17114 28314
rect 17166 28262 17178 28314
rect 17230 28262 17242 28314
rect 17294 28262 22922 28314
rect 22974 28262 22986 28314
rect 23038 28262 23050 28314
rect 23102 28262 23114 28314
rect 23166 28262 23178 28314
rect 23230 28262 23242 28314
rect 23294 28262 28922 28314
rect 28974 28262 28986 28314
rect 29038 28262 29050 28314
rect 29102 28262 29114 28314
rect 29166 28262 29178 28314
rect 29230 28262 29242 28314
rect 29294 28262 31832 28314
rect 1104 28240 31832 28262
rect 8478 28160 8484 28212
rect 8536 28200 8542 28212
rect 8757 28203 8815 28209
rect 8757 28200 8769 28203
rect 8536 28172 8769 28200
rect 8536 28160 8542 28172
rect 8757 28169 8769 28172
rect 8803 28169 8815 28203
rect 8757 28163 8815 28169
rect 10502 28160 10508 28212
rect 10560 28160 10566 28212
rect 13722 28160 13728 28212
rect 13780 28160 13786 28212
rect 13814 28160 13820 28212
rect 13872 28160 13878 28212
rect 14090 28160 14096 28212
rect 14148 28160 14154 28212
rect 14366 28160 14372 28212
rect 14424 28160 14430 28212
rect 14458 28160 14464 28212
rect 14516 28200 14522 28212
rect 14921 28203 14979 28209
rect 14921 28200 14933 28203
rect 14516 28172 14933 28200
rect 14516 28160 14522 28172
rect 14921 28169 14933 28172
rect 14967 28169 14979 28203
rect 14921 28163 14979 28169
rect 15028 28172 17908 28200
rect 9125 28067 9183 28073
rect 9125 28033 9137 28067
rect 9171 28064 9183 28067
rect 9769 28067 9827 28073
rect 9769 28064 9781 28067
rect 9171 28036 9781 28064
rect 9171 28033 9183 28036
rect 9125 28027 9183 28033
rect 9769 28033 9781 28036
rect 9815 28033 9827 28067
rect 9769 28027 9827 28033
rect 9214 27956 9220 28008
rect 9272 27956 9278 28008
rect 9309 27999 9367 28005
rect 9309 27965 9321 27999
rect 9355 27965 9367 27999
rect 9309 27959 9367 27965
rect 9324 27928 9352 27959
rect 9858 27956 9864 28008
rect 9916 27996 9922 28008
rect 10318 27996 10324 28008
rect 9916 27968 10324 27996
rect 9916 27956 9922 27968
rect 10318 27956 10324 27968
rect 10376 27956 10382 28008
rect 10520 28005 10548 28160
rect 14108 28132 14136 28160
rect 13372 28104 14136 28132
rect 14384 28132 14412 28160
rect 14829 28135 14887 28141
rect 14829 28132 14841 28135
rect 14384 28104 14841 28132
rect 10873 28067 10931 28073
rect 10873 28033 10885 28067
rect 10919 28064 10931 28067
rect 11609 28067 11667 28073
rect 11609 28064 11621 28067
rect 10919 28036 11621 28064
rect 10919 28033 10931 28036
rect 10873 28027 10931 28033
rect 11609 28033 11621 28036
rect 11655 28033 11667 28067
rect 11609 28027 11667 28033
rect 11882 28024 11888 28076
rect 11940 28064 11946 28076
rect 13372 28073 13400 28104
rect 14829 28101 14841 28104
rect 14875 28101 14887 28135
rect 14829 28095 14887 28101
rect 12161 28067 12219 28073
rect 12161 28064 12173 28067
rect 11940 28036 12173 28064
rect 11940 28024 11946 28036
rect 12161 28033 12173 28036
rect 12207 28033 12219 28067
rect 12161 28027 12219 28033
rect 13357 28067 13415 28073
rect 13357 28033 13369 28067
rect 13403 28033 13415 28067
rect 13357 28027 13415 28033
rect 13633 28067 13691 28073
rect 13633 28033 13645 28067
rect 13679 28064 13691 28067
rect 13906 28064 13912 28076
rect 13679 28036 13912 28064
rect 13679 28033 13691 28036
rect 13633 28027 13691 28033
rect 13906 28024 13912 28036
rect 13964 28024 13970 28076
rect 14274 28024 14280 28076
rect 14332 28024 14338 28076
rect 14366 28024 14372 28076
rect 14424 28024 14430 28076
rect 14461 28067 14519 28073
rect 14461 28033 14473 28067
rect 14507 28064 14519 28067
rect 14642 28064 14648 28076
rect 14507 28036 14648 28064
rect 14507 28033 14519 28036
rect 14461 28027 14519 28033
rect 14642 28024 14648 28036
rect 14700 28024 14706 28076
rect 10505 27999 10563 28005
rect 10505 27965 10517 27999
rect 10551 27965 10563 27999
rect 10505 27959 10563 27965
rect 10686 27956 10692 28008
rect 10744 27996 10750 28008
rect 10781 27999 10839 28005
rect 10781 27996 10793 27999
rect 10744 27968 10793 27996
rect 10744 27956 10750 27968
rect 10781 27965 10793 27968
rect 10827 27965 10839 27999
rect 13173 27999 13231 28005
rect 13173 27996 13185 27999
rect 10781 27959 10839 27965
rect 12406 27968 13185 27996
rect 12406 27928 12434 27968
rect 13173 27965 13185 27968
rect 13219 27996 13231 27999
rect 13722 27996 13728 28008
rect 13219 27968 13728 27996
rect 13219 27965 13231 27968
rect 13173 27959 13231 27965
rect 13722 27956 13728 27968
rect 13780 27956 13786 28008
rect 14734 27996 14740 28008
rect 14660 27968 14740 27996
rect 9232 27900 12434 27928
rect 7834 27820 7840 27872
rect 7892 27860 7898 27872
rect 9232 27860 9260 27900
rect 13998 27888 14004 27940
rect 14056 27928 14062 27940
rect 14366 27928 14372 27940
rect 14056 27900 14372 27928
rect 14056 27888 14062 27900
rect 14366 27888 14372 27900
rect 14424 27928 14430 27940
rect 14660 27937 14688 27968
rect 14734 27956 14740 27968
rect 14792 27996 14798 28008
rect 15028 27996 15056 28172
rect 16945 28135 17003 28141
rect 16945 28132 16957 28135
rect 16684 28104 16957 28132
rect 16684 28073 16712 28104
rect 16945 28101 16957 28104
rect 16991 28132 17003 28135
rect 17586 28132 17592 28144
rect 16991 28104 17592 28132
rect 16991 28101 17003 28104
rect 16945 28095 17003 28101
rect 17586 28092 17592 28104
rect 17644 28092 17650 28144
rect 17880 28073 17908 28172
rect 16669 28067 16727 28073
rect 16669 28064 16681 28067
rect 14792 27968 15056 27996
rect 16224 28036 16681 28064
rect 14792 27956 14798 27968
rect 16224 27937 16252 28036
rect 16669 28033 16681 28036
rect 16715 28033 16727 28067
rect 16669 28027 16727 28033
rect 16853 28067 16911 28073
rect 16853 28033 16865 28067
rect 16899 28033 16911 28067
rect 16853 28027 16911 28033
rect 17865 28067 17923 28073
rect 17865 28033 17877 28067
rect 17911 28064 17923 28067
rect 18874 28064 18880 28076
rect 17911 28036 18880 28064
rect 17911 28033 17923 28036
rect 17865 28027 17923 28033
rect 16485 27999 16543 28005
rect 16485 27965 16497 27999
rect 16531 27996 16543 27999
rect 16574 27996 16580 28008
rect 16531 27968 16580 27996
rect 16531 27965 16543 27968
rect 16485 27959 16543 27965
rect 16574 27956 16580 27968
rect 16632 27996 16638 28008
rect 16868 27996 16896 28027
rect 18874 28024 18880 28036
rect 18932 28024 18938 28076
rect 20346 28024 20352 28076
rect 20404 28024 20410 28076
rect 23382 28024 23388 28076
rect 23440 28024 23446 28076
rect 26602 28024 26608 28076
rect 26660 28024 26666 28076
rect 16632 27968 16896 27996
rect 16632 27956 16638 27968
rect 14645 27931 14703 27937
rect 14645 27928 14657 27931
rect 14424 27900 14657 27928
rect 14424 27888 14430 27900
rect 14645 27897 14657 27900
rect 14691 27897 14703 27931
rect 16209 27931 16267 27937
rect 14645 27891 14703 27897
rect 15212 27900 16160 27928
rect 7892 27832 9260 27860
rect 7892 27820 7898 27832
rect 11330 27820 11336 27872
rect 11388 27860 11394 27872
rect 13449 27863 13507 27869
rect 13449 27860 13461 27863
rect 11388 27832 13461 27860
rect 11388 27820 11394 27832
rect 13449 27829 13461 27832
rect 13495 27829 13507 27863
rect 13449 27823 13507 27829
rect 14090 27820 14096 27872
rect 14148 27820 14154 27872
rect 14274 27820 14280 27872
rect 14332 27860 14338 27872
rect 15212 27860 15240 27900
rect 14332 27832 15240 27860
rect 14332 27820 14338 27832
rect 15838 27820 15844 27872
rect 15896 27860 15902 27872
rect 16025 27863 16083 27869
rect 16025 27860 16037 27863
rect 15896 27832 16037 27860
rect 15896 27820 15902 27832
rect 16025 27829 16037 27832
rect 16071 27829 16083 27863
rect 16132 27860 16160 27900
rect 16209 27897 16221 27931
rect 16255 27897 16267 27931
rect 16868 27928 16896 27968
rect 16942 27956 16948 28008
rect 17000 27996 17006 28008
rect 17678 27996 17684 28008
rect 17000 27968 17684 27996
rect 17000 27956 17006 27968
rect 17678 27956 17684 27968
rect 17736 27956 17742 28008
rect 18046 27956 18052 28008
rect 18104 27996 18110 28008
rect 18966 27996 18972 28008
rect 18104 27968 18972 27996
rect 18104 27956 18110 27968
rect 18966 27956 18972 27968
rect 19024 27996 19030 28008
rect 20162 27996 20168 28008
rect 19024 27968 20168 27996
rect 19024 27956 19030 27968
rect 20162 27956 20168 27968
rect 20220 27996 20226 28008
rect 20257 27999 20315 28005
rect 20257 27996 20269 27999
rect 20220 27968 20269 27996
rect 20220 27956 20226 27968
rect 20257 27965 20269 27968
rect 20303 27965 20315 27999
rect 20257 27959 20315 27965
rect 17313 27931 17371 27937
rect 17313 27928 17325 27931
rect 16868 27900 17325 27928
rect 16209 27891 16267 27897
rect 17313 27897 17325 27900
rect 17359 27928 17371 27931
rect 19978 27928 19984 27940
rect 17359 27900 19984 27928
rect 17359 27897 17371 27900
rect 17313 27891 17371 27897
rect 19978 27888 19984 27900
rect 20036 27888 20042 27940
rect 20714 27888 20720 27940
rect 20772 27888 20778 27940
rect 16666 27860 16672 27872
rect 16132 27832 16672 27860
rect 16025 27823 16083 27829
rect 16666 27820 16672 27832
rect 16724 27820 16730 27872
rect 16758 27820 16764 27872
rect 16816 27860 16822 27872
rect 17405 27863 17463 27869
rect 17405 27860 17417 27863
rect 16816 27832 17417 27860
rect 16816 27820 16822 27832
rect 17405 27829 17417 27832
rect 17451 27829 17463 27863
rect 17405 27823 17463 27829
rect 17681 27863 17739 27869
rect 17681 27829 17693 27863
rect 17727 27860 17739 27863
rect 17770 27860 17776 27872
rect 17727 27832 17776 27860
rect 17727 27829 17739 27832
rect 17681 27823 17739 27829
rect 17770 27820 17776 27832
rect 17828 27820 17834 27872
rect 23106 27820 23112 27872
rect 23164 27860 23170 27872
rect 23201 27863 23259 27869
rect 23201 27860 23213 27863
rect 23164 27832 23213 27860
rect 23164 27820 23170 27832
rect 23201 27829 23213 27832
rect 23247 27829 23259 27863
rect 23201 27823 23259 27829
rect 26326 27820 26332 27872
rect 26384 27860 26390 27872
rect 26421 27863 26479 27869
rect 26421 27860 26433 27863
rect 26384 27832 26433 27860
rect 26384 27820 26390 27832
rect 26421 27829 26433 27832
rect 26467 27829 26479 27863
rect 26421 27823 26479 27829
rect 1104 27770 31832 27792
rect 1104 27718 4182 27770
rect 4234 27718 4246 27770
rect 4298 27718 4310 27770
rect 4362 27718 4374 27770
rect 4426 27718 4438 27770
rect 4490 27718 4502 27770
rect 4554 27718 10182 27770
rect 10234 27718 10246 27770
rect 10298 27718 10310 27770
rect 10362 27718 10374 27770
rect 10426 27718 10438 27770
rect 10490 27718 10502 27770
rect 10554 27718 16182 27770
rect 16234 27718 16246 27770
rect 16298 27718 16310 27770
rect 16362 27718 16374 27770
rect 16426 27718 16438 27770
rect 16490 27718 16502 27770
rect 16554 27718 22182 27770
rect 22234 27718 22246 27770
rect 22298 27718 22310 27770
rect 22362 27718 22374 27770
rect 22426 27718 22438 27770
rect 22490 27718 22502 27770
rect 22554 27718 28182 27770
rect 28234 27718 28246 27770
rect 28298 27718 28310 27770
rect 28362 27718 28374 27770
rect 28426 27718 28438 27770
rect 28490 27718 28502 27770
rect 28554 27718 31832 27770
rect 1104 27696 31832 27718
rect 14918 27616 14924 27668
rect 14976 27656 14982 27668
rect 15562 27656 15568 27668
rect 14976 27628 15568 27656
rect 14976 27616 14982 27628
rect 15562 27616 15568 27628
rect 15620 27656 15626 27668
rect 16482 27656 16488 27668
rect 15620 27628 16488 27656
rect 15620 27616 15626 27628
rect 16482 27616 16488 27628
rect 16540 27616 16546 27668
rect 16592 27628 17816 27656
rect 13924 27560 14755 27588
rect 13924 27532 13952 27560
rect 13906 27480 13912 27532
rect 13964 27480 13970 27532
rect 8662 27412 8668 27464
rect 8720 27452 8726 27464
rect 9033 27455 9091 27461
rect 9033 27452 9045 27455
rect 8720 27424 9045 27452
rect 8720 27412 8726 27424
rect 9033 27421 9045 27424
rect 9079 27421 9091 27455
rect 11057 27455 11115 27461
rect 11057 27452 11069 27455
rect 9033 27415 9091 27421
rect 10428 27424 11069 27452
rect 4798 27344 4804 27396
rect 4856 27384 4862 27396
rect 7101 27387 7159 27393
rect 7101 27384 7113 27387
rect 4856 27356 7113 27384
rect 4856 27344 4862 27356
rect 7101 27353 7113 27356
rect 7147 27353 7159 27387
rect 7101 27347 7159 27353
rect 7469 27387 7527 27393
rect 7469 27353 7481 27387
rect 7515 27384 7527 27387
rect 9122 27384 9128 27396
rect 7515 27356 9128 27384
rect 7515 27353 7527 27356
rect 7469 27347 7527 27353
rect 9122 27344 9128 27356
rect 9180 27344 9186 27396
rect 9306 27393 9312 27396
rect 9300 27347 9312 27393
rect 9306 27344 9312 27347
rect 9364 27344 9370 27396
rect 10042 27276 10048 27328
rect 10100 27316 10106 27328
rect 10428 27325 10456 27424
rect 11057 27421 11069 27424
rect 11103 27421 11115 27455
rect 11057 27415 11115 27421
rect 13817 27455 13875 27461
rect 13817 27421 13829 27455
rect 13863 27452 13875 27455
rect 14090 27452 14096 27464
rect 13863 27424 14096 27452
rect 13863 27421 13875 27424
rect 13817 27415 13875 27421
rect 14090 27412 14096 27424
rect 14148 27412 14154 27464
rect 10594 27344 10600 27396
rect 10652 27384 10658 27396
rect 13449 27387 13507 27393
rect 13449 27384 13461 27387
rect 10652 27356 13461 27384
rect 10652 27344 10658 27356
rect 13449 27353 13461 27356
rect 13495 27353 13507 27387
rect 14384 27384 14412 27560
rect 14458 27480 14464 27532
rect 14516 27480 14522 27532
rect 14727 27529 14755 27560
rect 15010 27548 15016 27600
rect 15068 27588 15074 27600
rect 16592 27588 16620 27628
rect 15068 27560 16620 27588
rect 15068 27548 15074 27560
rect 16666 27548 16672 27600
rect 16724 27588 16730 27600
rect 16761 27591 16819 27597
rect 16761 27588 16773 27591
rect 16724 27560 16773 27588
rect 16724 27548 16730 27560
rect 16761 27557 16773 27560
rect 16807 27557 16819 27591
rect 16761 27551 16819 27557
rect 16942 27548 16948 27600
rect 17000 27588 17006 27600
rect 17402 27588 17408 27600
rect 17000 27560 17408 27588
rect 17000 27548 17006 27560
rect 17402 27548 17408 27560
rect 17460 27548 17466 27600
rect 17788 27588 17816 27628
rect 17862 27616 17868 27668
rect 17920 27656 17926 27668
rect 18414 27656 18420 27668
rect 17920 27628 18420 27656
rect 17920 27616 17926 27628
rect 18414 27616 18420 27628
rect 18472 27616 18478 27668
rect 17788 27560 17908 27588
rect 14712 27523 14770 27529
rect 14712 27489 14724 27523
rect 14758 27489 14770 27523
rect 14712 27483 14770 27489
rect 16022 27480 16028 27532
rect 16080 27480 16086 27532
rect 17880 27520 17908 27560
rect 18322 27548 18328 27600
rect 18380 27588 18386 27600
rect 19702 27588 19708 27600
rect 18380 27560 19708 27588
rect 18380 27548 18386 27560
rect 19702 27548 19708 27560
rect 19760 27548 19766 27600
rect 19797 27591 19855 27597
rect 19797 27557 19809 27591
rect 19843 27588 19855 27591
rect 20717 27591 20775 27597
rect 20717 27588 20729 27591
rect 19843 27560 20729 27588
rect 19843 27557 19855 27560
rect 19797 27551 19855 27557
rect 20717 27557 20729 27560
rect 20763 27557 20775 27591
rect 20717 27551 20775 27557
rect 29362 27548 29368 27600
rect 29420 27588 29426 27600
rect 30558 27588 30564 27600
rect 29420 27560 30564 27588
rect 29420 27548 29426 27560
rect 30558 27548 30564 27560
rect 30616 27548 30622 27600
rect 16500 27492 17816 27520
rect 17880 27492 18828 27520
rect 14476 27452 14504 27480
rect 14921 27455 14979 27461
rect 14921 27452 14933 27455
rect 14476 27424 14933 27452
rect 14921 27421 14933 27424
rect 14967 27452 14979 27455
rect 15010 27452 15016 27464
rect 14967 27424 15016 27452
rect 14967 27421 14979 27424
rect 14921 27415 14979 27421
rect 15010 27412 15016 27424
rect 15068 27412 15074 27464
rect 15197 27455 15255 27461
rect 15197 27421 15209 27455
rect 15243 27452 15255 27455
rect 16040 27452 16068 27480
rect 16117 27455 16175 27461
rect 16117 27452 16129 27455
rect 15243 27424 16129 27452
rect 15243 27421 15255 27424
rect 15197 27415 15255 27421
rect 16117 27421 16129 27424
rect 16163 27421 16175 27455
rect 16117 27415 16175 27421
rect 16500 27384 16528 27492
rect 17788 27461 17816 27492
rect 16602 27455 16660 27461
rect 16602 27421 16614 27455
rect 16648 27452 16660 27455
rect 17773 27455 17831 27461
rect 16648 27424 17448 27452
rect 16648 27421 16660 27424
rect 16602 27415 16660 27421
rect 17420 27396 17448 27424
rect 17773 27421 17785 27455
rect 17819 27452 17831 27455
rect 17862 27452 17868 27464
rect 17819 27424 17868 27452
rect 17819 27421 17831 27424
rect 17773 27415 17831 27421
rect 17862 27412 17868 27424
rect 17920 27412 17926 27464
rect 18046 27412 18052 27464
rect 18104 27412 18110 27464
rect 18156 27424 18460 27452
rect 16758 27384 16764 27396
rect 14384 27356 16764 27384
rect 13449 27347 13507 27353
rect 16758 27344 16764 27356
rect 16816 27344 16822 27396
rect 17402 27344 17408 27396
rect 17460 27384 17466 27396
rect 17681 27387 17739 27393
rect 17681 27384 17693 27387
rect 17460 27356 17693 27384
rect 17460 27344 17466 27356
rect 17681 27353 17693 27356
rect 17727 27384 17739 27387
rect 18156 27384 18184 27424
rect 17727 27356 18184 27384
rect 17727 27353 17739 27356
rect 17681 27347 17739 27353
rect 18322 27344 18328 27396
rect 18380 27344 18386 27396
rect 18432 27384 18460 27424
rect 18506 27412 18512 27464
rect 18564 27452 18570 27464
rect 18693 27455 18751 27461
rect 18693 27452 18705 27455
rect 18564 27424 18705 27452
rect 18564 27412 18570 27424
rect 18693 27421 18705 27424
rect 18739 27421 18751 27455
rect 18693 27415 18751 27421
rect 18800 27384 18828 27492
rect 19334 27480 19340 27532
rect 19392 27480 19398 27532
rect 19978 27480 19984 27532
rect 20036 27480 20042 27532
rect 18966 27412 18972 27464
rect 19024 27412 19030 27464
rect 19429 27455 19487 27461
rect 19429 27421 19441 27455
rect 19475 27452 19487 27455
rect 19886 27452 19892 27464
rect 19475 27424 19892 27452
rect 19475 27421 19487 27424
rect 19429 27415 19487 27421
rect 19886 27412 19892 27424
rect 19944 27412 19950 27464
rect 20070 27412 20076 27464
rect 20128 27412 20134 27464
rect 20714 27412 20720 27464
rect 20772 27452 20778 27464
rect 20993 27455 21051 27461
rect 20993 27452 21005 27455
rect 20772 27424 21005 27452
rect 20772 27412 20778 27424
rect 20993 27421 21005 27424
rect 21039 27421 21051 27455
rect 20993 27415 21051 27421
rect 22830 27412 22836 27464
rect 22888 27412 22894 27464
rect 23106 27461 23112 27464
rect 23100 27452 23112 27461
rect 23067 27424 23112 27452
rect 23100 27415 23112 27424
rect 23106 27412 23112 27415
rect 23164 27412 23170 27464
rect 24949 27455 25007 27461
rect 24949 27452 24961 27455
rect 24228 27424 24961 27452
rect 21269 27387 21327 27393
rect 21269 27384 21281 27387
rect 18432 27356 18736 27384
rect 18800 27356 21281 27384
rect 18708 27328 18736 27356
rect 21269 27353 21281 27356
rect 21315 27353 21327 27387
rect 21269 27347 21327 27353
rect 24228 27328 24256 27424
rect 24949 27421 24961 27424
rect 24995 27421 25007 27455
rect 24949 27415 25007 27421
rect 25314 27412 25320 27464
rect 25372 27452 25378 27464
rect 26326 27461 26332 27464
rect 26053 27455 26111 27461
rect 26053 27452 26065 27455
rect 25372 27424 26065 27452
rect 25372 27412 25378 27424
rect 26053 27421 26065 27424
rect 26099 27421 26111 27455
rect 26320 27452 26332 27461
rect 26287 27424 26332 27452
rect 26053 27415 26111 27421
rect 26320 27415 26332 27424
rect 26326 27412 26332 27415
rect 26384 27412 26390 27464
rect 28077 27455 28135 27461
rect 28077 27452 28089 27455
rect 27448 27424 28089 27452
rect 10413 27319 10471 27325
rect 10413 27316 10425 27319
rect 10100 27288 10425 27316
rect 10100 27276 10106 27288
rect 10413 27285 10425 27288
rect 10459 27285 10471 27319
rect 10413 27279 10471 27285
rect 10502 27276 10508 27328
rect 10560 27276 10566 27328
rect 14550 27276 14556 27328
rect 14608 27276 14614 27328
rect 14829 27319 14887 27325
rect 14829 27285 14841 27319
rect 14875 27316 14887 27319
rect 15930 27316 15936 27328
rect 14875 27288 15936 27316
rect 14875 27285 14887 27288
rect 14829 27279 14887 27285
rect 15930 27276 15936 27288
rect 15988 27276 15994 27328
rect 16114 27276 16120 27328
rect 16172 27316 16178 27328
rect 16393 27319 16451 27325
rect 16393 27316 16405 27319
rect 16172 27288 16405 27316
rect 16172 27276 16178 27288
rect 16393 27285 16405 27288
rect 16439 27285 16451 27319
rect 16393 27279 16451 27285
rect 16482 27276 16488 27328
rect 16540 27276 16546 27328
rect 16574 27276 16580 27328
rect 16632 27316 16638 27328
rect 17589 27319 17647 27325
rect 17589 27316 17601 27319
rect 16632 27288 17601 27316
rect 16632 27276 16638 27288
rect 17589 27285 17601 27288
rect 17635 27285 17647 27319
rect 17589 27279 17647 27285
rect 17957 27319 18015 27325
rect 17957 27285 17969 27319
rect 18003 27316 18015 27319
rect 18598 27316 18604 27328
rect 18003 27288 18604 27316
rect 18003 27285 18015 27288
rect 17957 27279 18015 27285
rect 18598 27276 18604 27288
rect 18656 27276 18662 27328
rect 18690 27276 18696 27328
rect 18748 27276 18754 27328
rect 20441 27319 20499 27325
rect 20441 27285 20453 27319
rect 20487 27316 20499 27319
rect 20901 27319 20959 27325
rect 20901 27316 20913 27319
rect 20487 27288 20913 27316
rect 20487 27285 20499 27288
rect 20441 27279 20499 27285
rect 20901 27285 20913 27288
rect 20947 27285 20959 27319
rect 20901 27279 20959 27285
rect 21082 27276 21088 27328
rect 21140 27276 21146 27328
rect 24210 27276 24216 27328
rect 24268 27276 24274 27328
rect 24394 27276 24400 27328
rect 24452 27276 24458 27328
rect 27246 27276 27252 27328
rect 27304 27316 27310 27328
rect 27448 27325 27476 27424
rect 28077 27421 28089 27424
rect 28123 27421 28135 27455
rect 28077 27415 28135 27421
rect 27433 27319 27491 27325
rect 27433 27316 27445 27319
rect 27304 27288 27445 27316
rect 27304 27276 27310 27288
rect 27433 27285 27445 27288
rect 27479 27285 27491 27319
rect 27433 27279 27491 27285
rect 27522 27276 27528 27328
rect 27580 27276 27586 27328
rect 1104 27226 31832 27248
rect 1104 27174 4922 27226
rect 4974 27174 4986 27226
rect 5038 27174 5050 27226
rect 5102 27174 5114 27226
rect 5166 27174 5178 27226
rect 5230 27174 5242 27226
rect 5294 27174 10922 27226
rect 10974 27174 10986 27226
rect 11038 27174 11050 27226
rect 11102 27174 11114 27226
rect 11166 27174 11178 27226
rect 11230 27174 11242 27226
rect 11294 27174 16922 27226
rect 16974 27174 16986 27226
rect 17038 27174 17050 27226
rect 17102 27174 17114 27226
rect 17166 27174 17178 27226
rect 17230 27174 17242 27226
rect 17294 27174 22922 27226
rect 22974 27174 22986 27226
rect 23038 27174 23050 27226
rect 23102 27174 23114 27226
rect 23166 27174 23178 27226
rect 23230 27174 23242 27226
rect 23294 27174 28922 27226
rect 28974 27174 28986 27226
rect 29038 27174 29050 27226
rect 29102 27174 29114 27226
rect 29166 27174 29178 27226
rect 29230 27174 29242 27226
rect 29294 27174 31832 27226
rect 1104 27152 31832 27174
rect 9217 27115 9275 27121
rect 9217 27081 9229 27115
rect 9263 27112 9275 27115
rect 9306 27112 9312 27124
rect 9263 27084 9312 27112
rect 9263 27081 9275 27084
rect 9217 27075 9275 27081
rect 9306 27072 9312 27084
rect 9364 27072 9370 27124
rect 9861 27115 9919 27121
rect 9861 27081 9873 27115
rect 9907 27112 9919 27115
rect 10502 27112 10508 27124
rect 9907 27084 10508 27112
rect 9907 27081 9919 27084
rect 9861 27075 9919 27081
rect 10502 27072 10508 27084
rect 10560 27072 10566 27124
rect 15010 27072 15016 27124
rect 15068 27072 15074 27124
rect 17034 27112 17040 27124
rect 15856 27084 17040 27112
rect 15856 27056 15884 27084
rect 17034 27072 17040 27084
rect 17092 27072 17098 27124
rect 17221 27115 17279 27121
rect 17221 27081 17233 27115
rect 17267 27112 17279 27115
rect 18046 27112 18052 27124
rect 17267 27084 18052 27112
rect 17267 27081 17279 27084
rect 17221 27075 17279 27081
rect 18046 27072 18052 27084
rect 18104 27072 18110 27124
rect 18138 27072 18144 27124
rect 18196 27112 18202 27124
rect 18325 27115 18383 27121
rect 18325 27112 18337 27115
rect 18196 27084 18337 27112
rect 18196 27072 18202 27084
rect 18325 27081 18337 27084
rect 18371 27081 18383 27115
rect 18325 27075 18383 27081
rect 18417 27115 18475 27121
rect 18417 27081 18429 27115
rect 18463 27112 18475 27115
rect 18690 27112 18696 27124
rect 18463 27084 18696 27112
rect 18463 27081 18475 27084
rect 18417 27075 18475 27081
rect 18690 27072 18696 27084
rect 18748 27072 18754 27124
rect 20901 27115 20959 27121
rect 20901 27081 20913 27115
rect 20947 27112 20959 27115
rect 21082 27112 21088 27124
rect 20947 27084 21088 27112
rect 20947 27081 20959 27084
rect 20901 27075 20959 27081
rect 21082 27072 21088 27084
rect 21140 27072 21146 27124
rect 23293 27115 23351 27121
rect 23293 27081 23305 27115
rect 23339 27112 23351 27115
rect 23382 27112 23388 27124
rect 23339 27084 23388 27112
rect 23339 27081 23351 27084
rect 23293 27075 23351 27081
rect 23382 27072 23388 27084
rect 23440 27072 23446 27124
rect 23661 27115 23719 27121
rect 23661 27081 23673 27115
rect 23707 27112 23719 27115
rect 24394 27112 24400 27124
rect 23707 27084 24400 27112
rect 23707 27081 23719 27084
rect 23661 27075 23719 27081
rect 24394 27072 24400 27084
rect 24452 27072 24458 27124
rect 26602 27072 26608 27124
rect 26660 27112 26666 27124
rect 26973 27115 27031 27121
rect 26973 27112 26985 27115
rect 26660 27084 26985 27112
rect 26660 27072 26666 27084
rect 26973 27081 26985 27084
rect 27019 27081 27031 27115
rect 26973 27075 27031 27081
rect 27341 27115 27399 27121
rect 27341 27081 27353 27115
rect 27387 27112 27399 27115
rect 27522 27112 27528 27124
rect 27387 27084 27528 27112
rect 27387 27081 27399 27084
rect 27341 27075 27399 27081
rect 27522 27072 27528 27084
rect 27580 27072 27586 27124
rect 28537 27115 28595 27121
rect 28537 27081 28549 27115
rect 28583 27081 28595 27115
rect 29362 27112 29368 27124
rect 28537 27075 28595 27081
rect 28644 27084 29368 27112
rect 8113 27047 8171 27053
rect 8113 27013 8125 27047
rect 8159 27044 8171 27047
rect 11330 27044 11336 27056
rect 8159 27016 11336 27044
rect 8159 27013 8171 27016
rect 8113 27007 8171 27013
rect 11330 27004 11336 27016
rect 11388 27004 11394 27056
rect 13372 27016 14688 27044
rect 6086 26936 6092 26988
rect 6144 26976 6150 26988
rect 13372 26985 13400 27016
rect 7745 26979 7803 26985
rect 7745 26976 7757 26979
rect 6144 26948 7757 26976
rect 6144 26936 6150 26948
rect 7745 26945 7757 26948
rect 7791 26945 7803 26979
rect 7745 26939 7803 26945
rect 9401 26979 9459 26985
rect 9401 26945 9413 26979
rect 9447 26976 9459 26979
rect 13357 26979 13415 26985
rect 9447 26948 9536 26976
rect 9447 26945 9459 26948
rect 9401 26939 9459 26945
rect 7377 26911 7435 26917
rect 7377 26877 7389 26911
rect 7423 26908 7435 26911
rect 8386 26908 8392 26920
rect 7423 26880 8392 26908
rect 7423 26877 7435 26880
rect 7377 26871 7435 26877
rect 8386 26868 8392 26880
rect 8444 26868 8450 26920
rect 9508 26849 9536 26948
rect 13357 26945 13369 26979
rect 13403 26945 13415 26979
rect 13357 26939 13415 26945
rect 13630 26936 13636 26988
rect 13688 26976 13694 26988
rect 13725 26979 13783 26985
rect 13725 26976 13737 26979
rect 13688 26948 13737 26976
rect 13688 26936 13694 26948
rect 13725 26945 13737 26948
rect 13771 26976 13783 26979
rect 14369 26979 14427 26985
rect 14369 26976 14381 26979
rect 13771 26948 14381 26976
rect 13771 26945 13783 26948
rect 13725 26939 13783 26945
rect 14369 26945 14381 26948
rect 14415 26945 14427 26979
rect 14369 26939 14427 26945
rect 14660 26976 14688 27016
rect 14826 27004 14832 27056
rect 14884 27044 14890 27056
rect 15222 27047 15280 27053
rect 15222 27044 15234 27047
rect 14884 27016 15234 27044
rect 14884 27004 14890 27016
rect 15222 27013 15234 27016
rect 15268 27044 15280 27047
rect 15838 27044 15844 27056
rect 15268 27016 15844 27044
rect 15268 27013 15280 27016
rect 15222 27007 15280 27013
rect 15838 27004 15844 27016
rect 15896 27004 15902 27056
rect 15930 27004 15936 27056
rect 15988 27044 15994 27056
rect 16326 27047 16384 27053
rect 16326 27044 16338 27047
rect 15988 27016 16338 27044
rect 15988 27004 15994 27016
rect 16326 27013 16338 27016
rect 16372 27013 16384 27047
rect 16326 27007 16384 27013
rect 16669 27047 16727 27053
rect 16669 27013 16681 27047
rect 16715 27044 16727 27047
rect 16758 27044 16764 27056
rect 16715 27016 16764 27044
rect 16715 27013 16727 27016
rect 16669 27007 16727 27013
rect 16758 27004 16764 27016
rect 16816 27004 16822 27056
rect 17402 27044 17408 27056
rect 16960 27016 17408 27044
rect 14918 26976 14924 26988
rect 14660 26948 14924 26976
rect 9674 26868 9680 26920
rect 9732 26908 9738 26920
rect 9953 26911 10011 26917
rect 9953 26908 9965 26911
rect 9732 26880 9965 26908
rect 9732 26868 9738 26880
rect 9953 26877 9965 26880
rect 9999 26877 10011 26911
rect 9953 26871 10011 26877
rect 10137 26911 10195 26917
rect 10137 26877 10149 26911
rect 10183 26908 10195 26911
rect 10594 26908 10600 26920
rect 10183 26880 10600 26908
rect 10183 26877 10195 26880
rect 10137 26871 10195 26877
rect 10594 26868 10600 26880
rect 10652 26868 10658 26920
rect 12526 26868 12532 26920
rect 12584 26908 12590 26920
rect 13446 26908 13452 26920
rect 12584 26880 13452 26908
rect 12584 26868 12590 26880
rect 13446 26868 13452 26880
rect 13504 26908 13510 26920
rect 13909 26911 13967 26917
rect 13909 26908 13921 26911
rect 13504 26880 13921 26908
rect 13504 26868 13510 26880
rect 13909 26877 13921 26880
rect 13955 26877 13967 26911
rect 13909 26871 13967 26877
rect 14277 26911 14335 26917
rect 14277 26877 14289 26911
rect 14323 26908 14335 26911
rect 14660 26908 14688 26948
rect 14918 26936 14924 26948
rect 14976 26936 14982 26988
rect 15010 26936 15016 26988
rect 15068 26976 15074 26988
rect 16114 26976 16120 26988
rect 15068 26948 16120 26976
rect 15068 26936 15074 26948
rect 16114 26936 16120 26948
rect 16172 26936 16178 26988
rect 16574 26936 16580 26988
rect 16632 26976 16638 26988
rect 16960 26985 16988 27016
rect 17402 27004 17408 27016
rect 17460 27004 17466 27056
rect 17589 27047 17647 27053
rect 17589 27044 17601 27047
rect 17512 27016 17601 27044
rect 16853 26979 16911 26985
rect 16853 26976 16865 26979
rect 16632 26948 16865 26976
rect 16632 26936 16638 26948
rect 16853 26945 16865 26948
rect 16899 26945 16911 26979
rect 16853 26939 16911 26945
rect 16945 26979 17003 26985
rect 16945 26945 16957 26979
rect 16991 26945 17003 26979
rect 16945 26939 17003 26945
rect 17126 26936 17132 26988
rect 17184 26976 17190 26988
rect 17512 26976 17540 27016
rect 17589 27013 17601 27016
rect 17635 27013 17647 27047
rect 17589 27007 17647 27013
rect 18230 27004 18236 27056
rect 18288 27044 18294 27056
rect 19429 27047 19487 27053
rect 19429 27044 19441 27047
rect 18288 27016 19441 27044
rect 18288 27004 18294 27016
rect 19429 27013 19441 27016
rect 19475 27013 19487 27047
rect 25676 27047 25734 27053
rect 19429 27007 19487 27013
rect 23768 27016 25636 27044
rect 23768 26988 23796 27016
rect 17184 26948 17540 26976
rect 17184 26936 17190 26948
rect 17678 26936 17684 26988
rect 17736 26936 17742 26988
rect 17770 26936 17776 26988
rect 17828 26985 17834 26988
rect 17828 26979 17856 26985
rect 17844 26945 17856 26979
rect 17828 26939 17856 26945
rect 17828 26936 17834 26939
rect 18322 26936 18328 26988
rect 18380 26976 18386 26988
rect 18785 26979 18843 26985
rect 18785 26976 18797 26979
rect 18380 26948 18797 26976
rect 18380 26936 18386 26948
rect 18785 26945 18797 26948
rect 18831 26945 18843 26979
rect 18785 26939 18843 26945
rect 20530 26936 20536 26988
rect 20588 26936 20594 26988
rect 23750 26936 23756 26988
rect 23808 26936 23814 26988
rect 25608 26976 25636 27016
rect 25676 27013 25688 27047
rect 25722 27044 25734 27047
rect 28552 27044 28580 27075
rect 25722 27016 28580 27044
rect 25722 27013 25734 27016
rect 25676 27007 25734 27013
rect 27433 26979 27491 26985
rect 27433 26976 27445 26979
rect 25608 26948 27445 26976
rect 27433 26945 27445 26948
rect 27479 26976 27491 26979
rect 28644 26976 28672 27084
rect 29362 27072 29368 27084
rect 29420 27072 29426 27124
rect 27479 26948 28672 26976
rect 27479 26945 27491 26948
rect 27433 26939 27491 26945
rect 28718 26936 28724 26988
rect 28776 26936 28782 26988
rect 14323 26880 14688 26908
rect 14323 26877 14335 26880
rect 14277 26871 14335 26877
rect 14734 26868 14740 26920
rect 14792 26917 14798 26920
rect 14792 26911 14822 26917
rect 14810 26908 14822 26911
rect 14810 26880 15056 26908
rect 14810 26877 14822 26880
rect 14792 26871 14822 26877
rect 14792 26868 14798 26871
rect 9493 26843 9551 26849
rect 9493 26809 9505 26843
rect 9539 26809 9551 26843
rect 9493 26803 9551 26809
rect 12802 26800 12808 26852
rect 12860 26800 12866 26852
rect 15028 26840 15056 26880
rect 15102 26868 15108 26920
rect 15160 26868 15166 26920
rect 15841 26911 15899 26917
rect 15841 26877 15853 26911
rect 15887 26908 15899 26911
rect 16022 26908 16028 26920
rect 15887 26880 16028 26908
rect 15887 26877 15899 26880
rect 15841 26871 15899 26877
rect 15856 26840 15884 26871
rect 16022 26868 16028 26880
rect 16080 26868 16086 26920
rect 16209 26911 16267 26917
rect 16209 26877 16221 26911
rect 16255 26877 16267 26911
rect 16209 26871 16267 26877
rect 17313 26911 17371 26917
rect 17313 26877 17325 26911
rect 17359 26877 17371 26911
rect 18049 26911 18107 26917
rect 18049 26908 18061 26911
rect 17313 26871 17371 26877
rect 17880 26880 18061 26908
rect 15028 26812 15884 26840
rect 16224 26840 16252 26871
rect 16390 26840 16396 26852
rect 16224 26812 16396 26840
rect 6730 26732 6736 26784
rect 6788 26732 6794 26784
rect 14553 26775 14611 26781
rect 14553 26741 14565 26775
rect 14599 26772 14611 26775
rect 15010 26772 15016 26784
rect 14599 26744 15016 26772
rect 14599 26741 14611 26744
rect 14553 26735 14611 26741
rect 15010 26732 15016 26744
rect 15068 26732 15074 26784
rect 15378 26732 15384 26784
rect 15436 26732 15442 26784
rect 15856 26772 15884 26812
rect 16390 26800 16396 26812
rect 16448 26800 16454 26852
rect 16485 26843 16543 26849
rect 16485 26809 16497 26843
rect 16531 26840 16543 26843
rect 16850 26840 16856 26852
rect 16531 26812 16856 26840
rect 16531 26809 16543 26812
rect 16485 26803 16543 26809
rect 16850 26800 16856 26812
rect 16908 26800 16914 26852
rect 17328 26772 17356 26871
rect 17880 26772 17908 26880
rect 18049 26877 18061 26880
rect 18095 26877 18107 26911
rect 18049 26871 18107 26877
rect 18414 26868 18420 26920
rect 18472 26908 18478 26920
rect 18534 26911 18592 26917
rect 18534 26908 18546 26911
rect 18472 26880 18546 26908
rect 18472 26868 18478 26880
rect 18534 26877 18546 26880
rect 18580 26877 18592 26911
rect 18534 26871 18592 26877
rect 19061 26911 19119 26917
rect 19061 26877 19073 26911
rect 19107 26908 19119 26911
rect 19150 26908 19156 26920
rect 19107 26880 19156 26908
rect 19107 26877 19119 26880
rect 19061 26871 19119 26877
rect 19150 26868 19156 26880
rect 19208 26868 19214 26920
rect 20438 26868 20444 26920
rect 20496 26868 20502 26920
rect 23937 26911 23995 26917
rect 23937 26908 23949 26911
rect 22066 26880 23949 26908
rect 17957 26843 18015 26849
rect 17957 26809 17969 26843
rect 18003 26840 18015 26843
rect 19334 26840 19340 26852
rect 18003 26812 19340 26840
rect 18003 26809 18015 26812
rect 17957 26803 18015 26809
rect 19334 26800 19340 26812
rect 19392 26800 19398 26852
rect 22066 26840 22094 26880
rect 23937 26877 23949 26880
rect 23983 26908 23995 26911
rect 25222 26908 25228 26920
rect 23983 26880 25228 26908
rect 23983 26877 23995 26880
rect 23937 26871 23995 26877
rect 25222 26868 25228 26880
rect 25280 26868 25286 26920
rect 25314 26868 25320 26920
rect 25372 26908 25378 26920
rect 25409 26911 25467 26917
rect 25409 26908 25421 26911
rect 25372 26880 25421 26908
rect 25372 26868 25378 26880
rect 25409 26877 25421 26880
rect 25455 26877 25467 26911
rect 25409 26871 25467 26877
rect 27525 26911 27583 26917
rect 27525 26877 27537 26911
rect 27571 26908 27583 26911
rect 27706 26908 27712 26920
rect 27571 26880 27712 26908
rect 27571 26877 27583 26880
rect 27525 26871 27583 26877
rect 27706 26868 27712 26880
rect 27764 26868 27770 26920
rect 28353 26911 28411 26917
rect 28353 26877 28365 26911
rect 28399 26877 28411 26911
rect 28353 26871 28411 26877
rect 19628 26812 22094 26840
rect 26789 26843 26847 26849
rect 15856 26744 17908 26772
rect 18690 26732 18696 26784
rect 18748 26732 18754 26784
rect 18782 26732 18788 26784
rect 18840 26772 18846 26784
rect 19628 26772 19656 26812
rect 26789 26809 26801 26843
rect 26835 26840 26847 26843
rect 28368 26840 28396 26871
rect 26835 26812 28396 26840
rect 26835 26809 26847 26812
rect 26789 26803 26847 26809
rect 27540 26784 27568 26812
rect 18840 26744 19656 26772
rect 19705 26775 19763 26781
rect 18840 26732 18846 26744
rect 19705 26741 19717 26775
rect 19751 26772 19763 26775
rect 21174 26772 21180 26784
rect 19751 26744 21180 26772
rect 19751 26741 19763 26744
rect 19705 26735 19763 26741
rect 21174 26732 21180 26744
rect 21232 26732 21238 26784
rect 27522 26732 27528 26784
rect 27580 26732 27586 26784
rect 27798 26732 27804 26784
rect 27856 26732 27862 26784
rect 1104 26682 31832 26704
rect 1104 26630 4182 26682
rect 4234 26630 4246 26682
rect 4298 26630 4310 26682
rect 4362 26630 4374 26682
rect 4426 26630 4438 26682
rect 4490 26630 4502 26682
rect 4554 26630 10182 26682
rect 10234 26630 10246 26682
rect 10298 26630 10310 26682
rect 10362 26630 10374 26682
rect 10426 26630 10438 26682
rect 10490 26630 10502 26682
rect 10554 26630 16182 26682
rect 16234 26630 16246 26682
rect 16298 26630 16310 26682
rect 16362 26630 16374 26682
rect 16426 26630 16438 26682
rect 16490 26630 16502 26682
rect 16554 26630 22182 26682
rect 22234 26630 22246 26682
rect 22298 26630 22310 26682
rect 22362 26630 22374 26682
rect 22426 26630 22438 26682
rect 22490 26630 22502 26682
rect 22554 26630 28182 26682
rect 28234 26630 28246 26682
rect 28298 26630 28310 26682
rect 28362 26630 28374 26682
rect 28426 26630 28438 26682
rect 28490 26630 28502 26682
rect 28554 26630 31832 26682
rect 1104 26608 31832 26630
rect 6641 26571 6699 26577
rect 6641 26537 6653 26571
rect 6687 26568 6699 26571
rect 8386 26568 8392 26580
rect 6687 26540 8392 26568
rect 6687 26537 6699 26540
rect 6641 26531 6699 26537
rect 8386 26528 8392 26540
rect 8444 26528 8450 26580
rect 9122 26528 9128 26580
rect 9180 26568 9186 26580
rect 15289 26571 15347 26577
rect 15289 26568 15301 26571
rect 9180 26540 15301 26568
rect 9180 26528 9186 26540
rect 15289 26537 15301 26540
rect 15335 26537 15347 26571
rect 15289 26531 15347 26537
rect 18138 26528 18144 26580
rect 18196 26528 18202 26580
rect 18598 26528 18604 26580
rect 18656 26528 18662 26580
rect 18690 26528 18696 26580
rect 18748 26528 18754 26580
rect 19150 26528 19156 26580
rect 19208 26568 19214 26580
rect 27706 26568 27712 26580
rect 19208 26540 27712 26568
rect 19208 26528 19214 26540
rect 27706 26528 27712 26540
rect 27764 26528 27770 26580
rect 27798 26528 27804 26580
rect 27856 26528 27862 26580
rect 27985 26571 28043 26577
rect 27985 26537 27997 26571
rect 28031 26568 28043 26571
rect 28718 26568 28724 26580
rect 28031 26540 28724 26568
rect 28031 26537 28043 26540
rect 27985 26531 28043 26537
rect 28718 26528 28724 26540
rect 28776 26528 28782 26580
rect 8113 26503 8171 26509
rect 8113 26469 8125 26503
rect 8159 26469 8171 26503
rect 8113 26463 8171 26469
rect 8128 26432 8156 26463
rect 14550 26460 14556 26512
rect 14608 26460 14614 26512
rect 14918 26460 14924 26512
rect 14976 26460 14982 26512
rect 15841 26503 15899 26509
rect 15841 26469 15853 26503
rect 15887 26500 15899 26503
rect 16758 26500 16764 26512
rect 15887 26472 16764 26500
rect 15887 26469 15899 26472
rect 15841 26463 15899 26469
rect 16758 26460 16764 26472
rect 16816 26460 16822 26512
rect 17497 26503 17555 26509
rect 17497 26469 17509 26503
rect 17543 26500 17555 26503
rect 18230 26500 18236 26512
rect 17543 26472 18236 26500
rect 17543 26469 17555 26472
rect 17497 26463 17555 26469
rect 18230 26460 18236 26472
rect 18288 26460 18294 26512
rect 9493 26435 9551 26441
rect 9493 26432 9505 26435
rect 8128 26404 9505 26432
rect 9493 26401 9505 26404
rect 9539 26432 9551 26435
rect 9950 26432 9956 26444
rect 9539 26404 9956 26432
rect 9539 26401 9551 26404
rect 9493 26395 9551 26401
rect 9950 26392 9956 26404
rect 10008 26392 10014 26444
rect 14568 26432 14596 26460
rect 13372 26404 14596 26432
rect 5261 26367 5319 26373
rect 5261 26333 5273 26367
rect 5307 26364 5319 26367
rect 6733 26367 6791 26373
rect 6733 26364 6745 26367
rect 5307 26336 6745 26364
rect 5307 26333 5319 26336
rect 5261 26327 5319 26333
rect 6733 26333 6745 26336
rect 6779 26364 6791 26367
rect 7282 26364 7288 26376
rect 6779 26336 7288 26364
rect 6779 26333 6791 26336
rect 6733 26327 6791 26333
rect 5276 26296 5304 26327
rect 7282 26324 7288 26336
rect 7340 26324 7346 26376
rect 13372 26373 13400 26404
rect 14734 26392 14740 26444
rect 14792 26392 14798 26444
rect 14829 26435 14887 26441
rect 14829 26401 14841 26435
rect 14875 26432 14887 26435
rect 14936 26432 14964 26460
rect 14875 26404 14964 26432
rect 14875 26401 14887 26404
rect 14829 26395 14887 26401
rect 15102 26392 15108 26444
rect 15160 26392 15166 26444
rect 16022 26392 16028 26444
rect 16080 26432 16086 26444
rect 16853 26435 16911 26441
rect 16853 26432 16865 26435
rect 16080 26404 16865 26432
rect 16080 26392 16086 26404
rect 16853 26401 16865 26404
rect 16899 26401 16911 26435
rect 16853 26395 16911 26401
rect 17126 26392 17132 26444
rect 17184 26392 17190 26444
rect 17221 26435 17279 26441
rect 17221 26401 17233 26435
rect 17267 26432 17279 26435
rect 17770 26432 17776 26444
rect 17267 26404 17776 26432
rect 17267 26401 17279 26404
rect 17221 26395 17279 26401
rect 17770 26392 17776 26404
rect 17828 26392 17834 26444
rect 13357 26367 13415 26373
rect 13357 26333 13369 26367
rect 13403 26333 13415 26367
rect 13357 26327 13415 26333
rect 13906 26324 13912 26376
rect 13964 26324 13970 26376
rect 14274 26324 14280 26376
rect 14332 26324 14338 26376
rect 14553 26367 14611 26373
rect 14553 26333 14565 26367
rect 14599 26364 14611 26367
rect 14752 26364 14780 26392
rect 14599 26336 14780 26364
rect 14921 26367 14979 26373
rect 14599 26333 14611 26336
rect 14553 26327 14611 26333
rect 14921 26333 14933 26367
rect 14967 26364 14979 26367
rect 15120 26364 15148 26392
rect 17494 26364 17500 26376
rect 14967 26336 17500 26364
rect 14967 26333 14979 26336
rect 14921 26327 14979 26333
rect 4080 26268 5304 26296
rect 5528 26299 5586 26305
rect 3970 26188 3976 26240
rect 4028 26228 4034 26240
rect 4080 26228 4108 26268
rect 5528 26265 5540 26299
rect 5574 26296 5586 26299
rect 7000 26299 7058 26305
rect 5574 26268 6960 26296
rect 5574 26265 5586 26268
rect 5528 26259 5586 26265
rect 4028 26200 4108 26228
rect 6932 26228 6960 26268
rect 7000 26265 7012 26299
rect 7046 26296 7058 26299
rect 7098 26296 7104 26308
rect 7046 26268 7104 26296
rect 7046 26265 7058 26268
rect 7000 26259 7058 26265
rect 7098 26256 7104 26268
rect 7156 26256 7162 26308
rect 13081 26299 13139 26305
rect 13081 26296 13093 26299
rect 12406 26268 13093 26296
rect 7558 26228 7564 26240
rect 6932 26200 7564 26228
rect 4028 26188 4034 26200
rect 7558 26188 7564 26200
rect 7616 26188 7622 26240
rect 8570 26188 8576 26240
rect 8628 26228 8634 26240
rect 8941 26231 8999 26237
rect 8941 26228 8953 26231
rect 8628 26200 8953 26228
rect 8628 26188 8634 26200
rect 8941 26197 8953 26200
rect 8987 26197 8999 26231
rect 8941 26191 8999 26197
rect 11330 26188 11336 26240
rect 11388 26228 11394 26240
rect 12406 26228 12434 26268
rect 13081 26265 13093 26268
rect 13127 26265 13139 26299
rect 13081 26259 13139 26265
rect 13170 26256 13176 26308
rect 13228 26296 13234 26308
rect 13633 26299 13691 26305
rect 13633 26296 13645 26299
rect 13228 26268 13645 26296
rect 13228 26256 13234 26268
rect 13633 26265 13645 26268
rect 13679 26265 13691 26299
rect 14292 26296 14320 26324
rect 15488 26305 15516 26336
rect 17494 26324 17500 26336
rect 17552 26364 17558 26376
rect 17865 26367 17923 26373
rect 17865 26364 17877 26367
rect 17552 26336 17877 26364
rect 17552 26324 17558 26336
rect 17865 26333 17877 26336
rect 17911 26333 17923 26367
rect 17865 26327 17923 26333
rect 18046 26324 18052 26376
rect 18104 26364 18110 26376
rect 18233 26367 18291 26373
rect 18233 26364 18245 26367
rect 18104 26336 18245 26364
rect 18104 26324 18110 26336
rect 18233 26333 18245 26336
rect 18279 26333 18291 26367
rect 18233 26327 18291 26333
rect 15038 26299 15096 26305
rect 15038 26296 15050 26299
rect 14292 26268 15050 26296
rect 13633 26259 13691 26265
rect 15038 26265 15050 26268
rect 15084 26265 15096 26299
rect 15038 26259 15096 26265
rect 15473 26299 15531 26305
rect 15473 26265 15485 26299
rect 15519 26265 15531 26299
rect 15473 26259 15531 26265
rect 15562 26256 15568 26308
rect 15620 26256 15626 26308
rect 15657 26299 15715 26305
rect 15657 26265 15669 26299
rect 15703 26296 15715 26299
rect 15746 26296 15752 26308
rect 15703 26268 15752 26296
rect 15703 26265 15715 26268
rect 15657 26259 15715 26265
rect 15746 26256 15752 26268
rect 15804 26256 15810 26308
rect 17034 26256 17040 26308
rect 17092 26296 17098 26308
rect 17338 26299 17396 26305
rect 17338 26296 17350 26299
rect 17092 26268 17350 26296
rect 17092 26256 17098 26268
rect 17338 26265 17350 26268
rect 17384 26265 17396 26299
rect 17338 26259 17396 26265
rect 17586 26256 17592 26308
rect 17644 26256 17650 26308
rect 17678 26256 17684 26308
rect 17736 26296 17742 26308
rect 17957 26299 18015 26305
rect 17957 26296 17969 26299
rect 17736 26268 17969 26296
rect 17736 26256 17742 26268
rect 17957 26265 17969 26268
rect 18003 26265 18015 26299
rect 17957 26259 18015 26265
rect 18322 26256 18328 26308
rect 18380 26296 18386 26308
rect 18509 26299 18567 26305
rect 18509 26296 18521 26299
rect 18380 26268 18521 26296
rect 18380 26256 18386 26268
rect 18509 26265 18521 26268
rect 18555 26265 18567 26299
rect 18616 26296 18644 26528
rect 18708 26364 18736 26528
rect 24486 26432 24492 26444
rect 22066 26404 24492 26432
rect 19337 26367 19395 26373
rect 19337 26364 19349 26367
rect 18708 26336 19349 26364
rect 19337 26333 19349 26336
rect 19383 26333 19395 26367
rect 19337 26327 19395 26333
rect 19705 26367 19763 26373
rect 19705 26333 19717 26367
rect 19751 26364 19763 26367
rect 22066 26364 22094 26404
rect 24486 26392 24492 26404
rect 24544 26392 24550 26444
rect 25314 26392 25320 26444
rect 25372 26432 25378 26444
rect 25777 26435 25835 26441
rect 25777 26432 25789 26435
rect 25372 26404 25789 26432
rect 25372 26392 25378 26404
rect 25777 26401 25789 26404
rect 25823 26401 25835 26435
rect 25777 26395 25835 26401
rect 27430 26392 27436 26444
rect 27488 26392 27494 26444
rect 19751 26336 22094 26364
rect 19751 26333 19763 26336
rect 19705 26327 19763 26333
rect 23474 26324 23480 26376
rect 23532 26324 23538 26376
rect 23658 26324 23664 26376
rect 23716 26324 23722 26376
rect 24302 26324 24308 26376
rect 24360 26364 24366 26376
rect 24949 26367 25007 26373
rect 24949 26364 24961 26367
rect 24360 26336 24961 26364
rect 24360 26324 24366 26336
rect 24949 26333 24961 26336
rect 24995 26333 25007 26367
rect 27448 26364 27476 26392
rect 24949 26327 25007 26333
rect 25056 26336 27476 26364
rect 27617 26367 27675 26373
rect 19889 26299 19947 26305
rect 19889 26296 19901 26299
rect 18616 26268 19901 26296
rect 18509 26259 18567 26265
rect 19889 26265 19901 26268
rect 19935 26265 19947 26299
rect 20254 26296 20260 26308
rect 19889 26259 19947 26265
rect 19996 26268 20260 26296
rect 11388 26200 12434 26228
rect 11388 26188 11394 26200
rect 15194 26188 15200 26240
rect 15252 26188 15258 26240
rect 15764 26228 15792 26256
rect 16482 26228 16488 26240
rect 15764 26200 16488 26228
rect 16482 26188 16488 26200
rect 16540 26228 16546 26240
rect 17773 26231 17831 26237
rect 17773 26228 17785 26231
rect 16540 26200 17785 26228
rect 16540 26188 16546 26200
rect 17773 26197 17785 26200
rect 17819 26197 17831 26231
rect 18524 26228 18552 26259
rect 18782 26228 18788 26240
rect 18524 26200 18788 26228
rect 17773 26191 17831 26197
rect 18782 26188 18788 26200
rect 18840 26188 18846 26240
rect 19702 26188 19708 26240
rect 19760 26228 19766 26240
rect 19996 26228 20024 26268
rect 20254 26256 20260 26268
rect 20312 26296 20318 26308
rect 25056 26296 25084 26336
rect 27617 26333 27629 26367
rect 27663 26364 27675 26367
rect 27816 26364 27844 26528
rect 27663 26336 27844 26364
rect 27663 26333 27675 26336
rect 27617 26327 27675 26333
rect 20312 26268 25084 26296
rect 26044 26299 26102 26305
rect 20312 26256 20318 26268
rect 26044 26265 26056 26299
rect 26090 26296 26102 26299
rect 26142 26296 26148 26308
rect 26090 26268 26148 26296
rect 26090 26265 26102 26268
rect 26044 26259 26102 26265
rect 26142 26256 26148 26268
rect 26200 26256 26206 26308
rect 31110 26256 31116 26308
rect 31168 26256 31174 26308
rect 31478 26256 31484 26308
rect 31536 26256 31542 26308
rect 19760 26200 20024 26228
rect 19760 26188 19766 26200
rect 20162 26188 20168 26240
rect 20220 26188 20226 26240
rect 23293 26231 23351 26237
rect 23293 26197 23305 26231
rect 23339 26228 23351 26231
rect 23382 26228 23388 26240
rect 23339 26200 23388 26228
rect 23339 26197 23351 26200
rect 23293 26191 23351 26197
rect 23382 26188 23388 26200
rect 23440 26188 23446 26240
rect 23845 26231 23903 26237
rect 23845 26197 23857 26231
rect 23891 26228 23903 26231
rect 24026 26228 24032 26240
rect 23891 26200 24032 26228
rect 23891 26197 23903 26200
rect 23845 26191 23903 26197
rect 24026 26188 24032 26200
rect 24084 26188 24090 26240
rect 24394 26188 24400 26240
rect 24452 26188 24458 26240
rect 26878 26188 26884 26240
rect 26936 26228 26942 26240
rect 27157 26231 27215 26237
rect 27157 26228 27169 26231
rect 26936 26200 27169 26228
rect 26936 26188 26942 26200
rect 27157 26197 27169 26200
rect 27203 26197 27215 26231
rect 27157 26191 27215 26197
rect 27525 26231 27583 26237
rect 27525 26197 27537 26231
rect 27571 26228 27583 26231
rect 27706 26228 27712 26240
rect 27571 26200 27712 26228
rect 27571 26197 27583 26200
rect 27525 26191 27583 26197
rect 27706 26188 27712 26200
rect 27764 26188 27770 26240
rect 1104 26138 31832 26160
rect 1104 26086 4922 26138
rect 4974 26086 4986 26138
rect 5038 26086 5050 26138
rect 5102 26086 5114 26138
rect 5166 26086 5178 26138
rect 5230 26086 5242 26138
rect 5294 26086 10922 26138
rect 10974 26086 10986 26138
rect 11038 26086 11050 26138
rect 11102 26086 11114 26138
rect 11166 26086 11178 26138
rect 11230 26086 11242 26138
rect 11294 26086 16922 26138
rect 16974 26086 16986 26138
rect 17038 26086 17050 26138
rect 17102 26086 17114 26138
rect 17166 26086 17178 26138
rect 17230 26086 17242 26138
rect 17294 26086 22922 26138
rect 22974 26086 22986 26138
rect 23038 26086 23050 26138
rect 23102 26086 23114 26138
rect 23166 26086 23178 26138
rect 23230 26086 23242 26138
rect 23294 26086 28922 26138
rect 28974 26086 28986 26138
rect 29038 26086 29050 26138
rect 29102 26086 29114 26138
rect 29166 26086 29178 26138
rect 29230 26086 29242 26138
rect 29294 26086 31832 26138
rect 1104 26064 31832 26086
rect 6730 25984 6736 26036
rect 6788 25984 6794 26036
rect 7098 25984 7104 26036
rect 7156 26024 7162 26036
rect 7285 26027 7343 26033
rect 7285 26024 7297 26027
rect 7156 25996 7297 26024
rect 7156 25984 7162 25996
rect 7285 25993 7297 25996
rect 7331 25993 7343 26027
rect 7285 25987 7343 25993
rect 7558 25984 7564 26036
rect 7616 25984 7622 26036
rect 7837 26027 7895 26033
rect 7837 25993 7849 26027
rect 7883 25993 7895 26027
rect 7837 25987 7895 25993
rect 8205 26027 8263 26033
rect 8205 25993 8217 26027
rect 8251 26024 8263 26027
rect 8570 26024 8576 26036
rect 8251 25996 8576 26024
rect 8251 25993 8263 25996
rect 8205 25987 8263 25993
rect 4893 25959 4951 25965
rect 4893 25925 4905 25959
rect 4939 25956 4951 25959
rect 5902 25956 5908 25968
rect 4939 25928 5908 25956
rect 4939 25925 4951 25928
rect 4893 25919 4951 25925
rect 5902 25916 5908 25928
rect 5960 25956 5966 25968
rect 6641 25959 6699 25965
rect 6641 25956 6653 25959
rect 5960 25928 6653 25956
rect 5960 25916 5966 25928
rect 6641 25925 6653 25928
rect 6687 25925 6699 25959
rect 7852 25956 7880 25987
rect 8570 25984 8576 25996
rect 8628 25984 8634 26036
rect 13906 25984 13912 26036
rect 13964 26024 13970 26036
rect 14093 26027 14151 26033
rect 14093 26024 14105 26027
rect 13964 25996 14105 26024
rect 13964 25984 13970 25996
rect 14093 25993 14105 25996
rect 14139 25993 14151 26027
rect 14093 25987 14151 25993
rect 14277 26027 14335 26033
rect 14277 25993 14289 26027
rect 14323 26024 14335 26027
rect 14826 26024 14832 26036
rect 14323 25996 14832 26024
rect 14323 25993 14335 25996
rect 14277 25987 14335 25993
rect 14826 25984 14832 25996
rect 14884 25984 14890 26036
rect 14918 25984 14924 26036
rect 14976 25984 14982 26036
rect 16666 25984 16672 26036
rect 16724 26024 16730 26036
rect 18046 26024 18052 26036
rect 16724 25996 18052 26024
rect 16724 25984 16730 25996
rect 18046 25984 18052 25996
rect 18104 25984 18110 26036
rect 21174 25984 21180 26036
rect 21232 26024 21238 26036
rect 22002 26024 22008 26036
rect 21232 25996 22008 26024
rect 21232 25984 21238 25996
rect 22002 25984 22008 25996
rect 22060 26024 22066 26036
rect 25590 26024 25596 26036
rect 22060 25996 25596 26024
rect 22060 25984 22066 25996
rect 25590 25984 25596 25996
rect 25648 25984 25654 26036
rect 6641 25919 6699 25925
rect 7484 25928 7880 25956
rect 9953 25959 10011 25965
rect 7484 25897 7512 25928
rect 9953 25925 9965 25959
rect 9999 25956 10011 25959
rect 14369 25959 14427 25965
rect 9999 25928 10732 25956
rect 9999 25925 10011 25928
rect 9953 25919 10011 25925
rect 10704 25900 10732 25928
rect 14369 25925 14381 25959
rect 14415 25956 14427 25959
rect 14936 25956 14964 25984
rect 14415 25928 14964 25956
rect 15105 25959 15163 25965
rect 14415 25925 14427 25928
rect 14369 25919 14427 25925
rect 15105 25925 15117 25959
rect 15151 25956 15163 25959
rect 15194 25956 15200 25968
rect 15151 25928 15200 25956
rect 15151 25925 15163 25928
rect 15105 25919 15163 25925
rect 15194 25916 15200 25928
rect 15252 25916 15258 25968
rect 15378 25916 15384 25968
rect 15436 25916 15442 25968
rect 19334 25916 19340 25968
rect 19392 25956 19398 25968
rect 19521 25959 19579 25965
rect 19521 25956 19533 25959
rect 19392 25928 19533 25956
rect 19392 25916 19398 25928
rect 19521 25925 19533 25928
rect 19567 25925 19579 25959
rect 25314 25956 25320 25968
rect 19521 25919 19579 25925
rect 23032 25928 25320 25956
rect 4525 25891 4583 25897
rect 4525 25857 4537 25891
rect 4571 25857 4583 25891
rect 4525 25851 4583 25857
rect 4985 25891 5043 25897
rect 4985 25857 4997 25891
rect 5031 25888 5043 25891
rect 5445 25891 5503 25897
rect 5445 25888 5457 25891
rect 5031 25860 5457 25888
rect 5031 25857 5043 25860
rect 4985 25851 5043 25857
rect 5445 25857 5457 25860
rect 5491 25857 5503 25891
rect 5445 25851 5503 25857
rect 7469 25891 7527 25897
rect 7469 25857 7481 25891
rect 7515 25857 7527 25891
rect 7469 25851 7527 25857
rect 7745 25891 7803 25897
rect 7745 25857 7757 25891
rect 7791 25857 7803 25891
rect 7745 25851 7803 25857
rect 4540 25752 4568 25851
rect 4798 25780 4804 25832
rect 4856 25780 4862 25832
rect 5994 25780 6000 25832
rect 6052 25780 6058 25832
rect 6549 25823 6607 25829
rect 6549 25789 6561 25823
rect 6595 25789 6607 25823
rect 7760 25820 7788 25851
rect 9674 25848 9680 25900
rect 9732 25848 9738 25900
rect 9858 25897 9864 25900
rect 9825 25891 9864 25897
rect 9825 25857 9837 25891
rect 9825 25851 9864 25857
rect 9858 25848 9864 25851
rect 9916 25848 9922 25900
rect 10042 25848 10048 25900
rect 10100 25848 10106 25900
rect 10134 25848 10140 25900
rect 10192 25897 10198 25900
rect 10192 25888 10200 25897
rect 10192 25860 10237 25888
rect 10192 25851 10200 25860
rect 10192 25848 10198 25851
rect 10686 25848 10692 25900
rect 10744 25848 10750 25900
rect 14461 25891 14519 25897
rect 14461 25857 14473 25891
rect 14507 25888 14519 25891
rect 14642 25888 14648 25900
rect 14507 25860 14648 25888
rect 14507 25857 14519 25860
rect 14461 25851 14519 25857
rect 14642 25848 14648 25860
rect 14700 25848 14706 25900
rect 18230 25848 18236 25900
rect 18288 25888 18294 25900
rect 18877 25891 18935 25897
rect 18877 25888 18889 25891
rect 18288 25860 18889 25888
rect 18288 25848 18294 25860
rect 18877 25857 18889 25860
rect 18923 25857 18935 25891
rect 18877 25851 18935 25857
rect 22830 25848 22836 25900
rect 22888 25848 22894 25900
rect 6549 25783 6607 25789
rect 7116 25792 7788 25820
rect 5442 25752 5448 25764
rect 4540 25724 5448 25752
rect 5442 25712 5448 25724
rect 5500 25712 5506 25764
rect 6564 25752 6592 25783
rect 7116 25761 7144 25792
rect 8294 25780 8300 25832
rect 8352 25780 8358 25832
rect 8481 25823 8539 25829
rect 8481 25789 8493 25823
rect 8527 25820 8539 25823
rect 13170 25820 13176 25832
rect 8527 25792 13176 25820
rect 8527 25789 8539 25792
rect 8481 25783 8539 25789
rect 13170 25780 13176 25792
rect 13228 25780 13234 25832
rect 14366 25780 14372 25832
rect 14424 25780 14430 25832
rect 19153 25823 19211 25829
rect 19153 25789 19165 25823
rect 19199 25820 19211 25823
rect 22646 25820 22652 25832
rect 19199 25792 22652 25820
rect 19199 25789 19211 25792
rect 19153 25783 19211 25789
rect 22646 25780 22652 25792
rect 22704 25780 22710 25832
rect 22848 25820 22876 25848
rect 22925 25823 22983 25829
rect 22925 25820 22937 25823
rect 22848 25792 22937 25820
rect 22925 25789 22937 25792
rect 22971 25820 22983 25823
rect 23032 25820 23060 25928
rect 23198 25897 23204 25900
rect 23192 25851 23204 25897
rect 23198 25848 23204 25851
rect 23256 25848 23262 25900
rect 24412 25897 24440 25928
rect 25314 25916 25320 25928
rect 25372 25916 25378 25968
rect 28994 25956 29000 25968
rect 26206 25928 29000 25956
rect 24397 25891 24455 25897
rect 24397 25857 24409 25891
rect 24443 25857 24455 25891
rect 24653 25891 24711 25897
rect 24653 25888 24665 25891
rect 24397 25851 24455 25857
rect 24504 25860 24665 25888
rect 22971 25792 23060 25820
rect 22971 25789 22983 25792
rect 22925 25783 22983 25789
rect 24026 25780 24032 25832
rect 24084 25820 24090 25832
rect 24504 25820 24532 25860
rect 24653 25857 24665 25860
rect 24699 25857 24711 25891
rect 26206 25888 26234 25928
rect 28994 25916 29000 25928
rect 29052 25916 29058 25968
rect 29181 25959 29239 25965
rect 29181 25925 29193 25959
rect 29227 25956 29239 25959
rect 29362 25956 29368 25968
rect 29227 25928 29368 25956
rect 29227 25925 29239 25928
rect 29181 25919 29239 25925
rect 29362 25916 29368 25928
rect 29420 25916 29426 25968
rect 24653 25851 24711 25857
rect 25424 25860 26234 25888
rect 26421 25891 26479 25897
rect 24084 25792 24532 25820
rect 24084 25780 24090 25792
rect 7101 25755 7159 25761
rect 6564 25724 6914 25752
rect 4341 25687 4399 25693
rect 4341 25653 4353 25687
rect 4387 25684 4399 25687
rect 4614 25684 4620 25696
rect 4387 25656 4620 25684
rect 4387 25653 4399 25656
rect 4341 25647 4399 25653
rect 4614 25644 4620 25656
rect 4672 25644 4678 25696
rect 5353 25687 5411 25693
rect 5353 25653 5365 25687
rect 5399 25684 5411 25687
rect 5534 25684 5540 25696
rect 5399 25656 5540 25684
rect 5399 25653 5411 25656
rect 5353 25647 5411 25653
rect 5534 25644 5540 25656
rect 5592 25644 5598 25696
rect 6886 25684 6914 25724
rect 7101 25721 7113 25755
rect 7147 25721 7159 25755
rect 11330 25752 11336 25764
rect 7101 25715 7159 25721
rect 7208 25724 11336 25752
rect 7208 25684 7236 25724
rect 11330 25712 11336 25724
rect 11388 25752 11394 25764
rect 11606 25752 11612 25764
rect 11388 25724 11612 25752
rect 11388 25712 11394 25724
rect 11606 25712 11612 25724
rect 11664 25712 11670 25764
rect 14384 25752 14412 25780
rect 14645 25755 14703 25761
rect 14645 25752 14657 25755
rect 14384 25724 14657 25752
rect 14645 25721 14657 25724
rect 14691 25721 14703 25755
rect 14645 25715 14703 25721
rect 24302 25712 24308 25764
rect 24360 25712 24366 25764
rect 6886 25656 7236 25684
rect 9490 25644 9496 25696
rect 9548 25684 9554 25696
rect 10134 25684 10140 25696
rect 9548 25656 10140 25684
rect 9548 25644 9554 25656
rect 10134 25644 10140 25656
rect 10192 25644 10198 25696
rect 10321 25687 10379 25693
rect 10321 25653 10333 25687
rect 10367 25684 10379 25687
rect 11422 25684 11428 25696
rect 10367 25656 11428 25684
rect 10367 25653 10379 25656
rect 10321 25647 10379 25653
rect 11422 25644 11428 25656
rect 11480 25644 11486 25696
rect 12158 25644 12164 25696
rect 12216 25684 12222 25696
rect 14829 25687 14887 25693
rect 14829 25684 14841 25687
rect 12216 25656 14841 25684
rect 12216 25644 12222 25656
rect 14829 25653 14841 25656
rect 14875 25653 14887 25687
rect 14829 25647 14887 25653
rect 15654 25644 15660 25696
rect 15712 25644 15718 25696
rect 19797 25687 19855 25693
rect 19797 25653 19809 25687
rect 19843 25684 19855 25687
rect 25424 25684 25452 25860
rect 26421 25857 26433 25891
rect 26467 25888 26479 25891
rect 26973 25891 27031 25897
rect 26973 25888 26985 25891
rect 26467 25860 26985 25888
rect 26467 25857 26479 25860
rect 26421 25851 26479 25857
rect 26973 25857 26985 25860
rect 27019 25857 27031 25891
rect 26973 25851 27031 25857
rect 26513 25823 26571 25829
rect 26513 25820 26525 25823
rect 25516 25792 26525 25820
rect 25516 25696 25544 25792
rect 26513 25789 26525 25792
rect 26559 25789 26571 25823
rect 26513 25783 26571 25789
rect 26697 25823 26755 25829
rect 26697 25789 26709 25823
rect 26743 25820 26755 25823
rect 26786 25820 26792 25832
rect 26743 25792 26792 25820
rect 26743 25789 26755 25792
rect 26697 25783 26755 25789
rect 25590 25712 25596 25764
rect 25648 25752 25654 25764
rect 26528 25752 26556 25783
rect 26786 25780 26792 25792
rect 26844 25780 26850 25832
rect 26878 25780 26884 25832
rect 26936 25820 26942 25832
rect 27617 25823 27675 25829
rect 27617 25820 27629 25823
rect 26936 25792 27629 25820
rect 26936 25780 26942 25792
rect 27617 25789 27629 25792
rect 27663 25789 27675 25823
rect 27617 25783 27675 25789
rect 27706 25752 27712 25764
rect 25648 25724 26234 25752
rect 26528 25724 27712 25752
rect 25648 25712 25654 25724
rect 19843 25656 25452 25684
rect 19843 25653 19855 25656
rect 19797 25647 19855 25653
rect 25498 25644 25504 25696
rect 25556 25644 25562 25696
rect 25774 25644 25780 25696
rect 25832 25644 25838 25696
rect 26050 25644 26056 25696
rect 26108 25644 26114 25696
rect 26206 25684 26234 25724
rect 27706 25712 27712 25724
rect 27764 25752 27770 25764
rect 29362 25752 29368 25764
rect 27764 25724 29368 25752
rect 27764 25712 27770 25724
rect 29362 25712 29368 25724
rect 29420 25712 29426 25764
rect 26786 25684 26792 25696
rect 26206 25656 26792 25684
rect 26786 25644 26792 25656
rect 26844 25644 26850 25696
rect 1104 25594 31832 25616
rect 1104 25542 4182 25594
rect 4234 25542 4246 25594
rect 4298 25542 4310 25594
rect 4362 25542 4374 25594
rect 4426 25542 4438 25594
rect 4490 25542 4502 25594
rect 4554 25542 10182 25594
rect 10234 25542 10246 25594
rect 10298 25542 10310 25594
rect 10362 25542 10374 25594
rect 10426 25542 10438 25594
rect 10490 25542 10502 25594
rect 10554 25542 16182 25594
rect 16234 25542 16246 25594
rect 16298 25542 16310 25594
rect 16362 25542 16374 25594
rect 16426 25542 16438 25594
rect 16490 25542 16502 25594
rect 16554 25542 22182 25594
rect 22234 25542 22246 25594
rect 22298 25542 22310 25594
rect 22362 25542 22374 25594
rect 22426 25542 22438 25594
rect 22490 25542 22502 25594
rect 22554 25542 28182 25594
rect 28234 25542 28246 25594
rect 28298 25542 28310 25594
rect 28362 25542 28374 25594
rect 28426 25542 28438 25594
rect 28490 25542 28502 25594
rect 28554 25542 31832 25594
rect 1104 25520 31832 25542
rect 5442 25440 5448 25492
rect 5500 25440 5506 25492
rect 5994 25440 6000 25492
rect 6052 25440 6058 25492
rect 9214 25480 9220 25492
rect 6104 25452 9220 25480
rect 5353 25415 5411 25421
rect 5353 25381 5365 25415
rect 5399 25412 5411 25415
rect 5626 25412 5632 25424
rect 5399 25384 5632 25412
rect 5399 25381 5411 25384
rect 5353 25375 5411 25381
rect 5626 25372 5632 25384
rect 5684 25412 5690 25424
rect 6012 25412 6040 25440
rect 5684 25384 6040 25412
rect 5684 25372 5690 25384
rect 3970 25304 3976 25356
rect 4028 25304 4034 25356
rect 5902 25304 5908 25356
rect 5960 25304 5966 25356
rect 5994 25304 6000 25356
rect 6052 25304 6058 25356
rect 5920 25276 5948 25304
rect 6104 25276 6132 25452
rect 9214 25440 9220 25452
rect 9272 25440 9278 25492
rect 9674 25440 9680 25492
rect 9732 25440 9738 25492
rect 20162 25440 20168 25492
rect 20220 25480 20226 25492
rect 20220 25452 22109 25480
rect 20220 25440 20226 25452
rect 8386 25372 8392 25424
rect 8444 25372 8450 25424
rect 9858 25372 9864 25424
rect 9916 25412 9922 25424
rect 10686 25412 10692 25424
rect 9916 25384 10692 25412
rect 9916 25372 9922 25384
rect 10686 25372 10692 25384
rect 10744 25372 10750 25424
rect 12161 25415 12219 25421
rect 12161 25381 12173 25415
rect 12207 25381 12219 25415
rect 12161 25375 12219 25381
rect 8404 25344 8432 25372
rect 8404 25316 10272 25344
rect 5920 25248 6132 25276
rect 6914 25236 6920 25288
rect 6972 25236 6978 25288
rect 7282 25236 7288 25288
rect 7340 25276 7346 25288
rect 8662 25276 8668 25288
rect 7340 25248 8668 25276
rect 7340 25236 7346 25248
rect 8662 25236 8668 25248
rect 8720 25236 8726 25288
rect 9493 25279 9551 25285
rect 9493 25245 9505 25279
rect 9539 25245 9551 25279
rect 9861 25279 9919 25285
rect 9861 25276 9873 25279
rect 9493 25239 9551 25245
rect 9646 25248 9873 25276
rect 4240 25211 4298 25217
rect 4240 25177 4252 25211
rect 4286 25208 4298 25211
rect 4798 25208 4804 25220
rect 4286 25180 4804 25208
rect 4286 25177 4298 25180
rect 4240 25171 4298 25177
rect 4798 25168 4804 25180
rect 4856 25168 4862 25220
rect 5813 25211 5871 25217
rect 5813 25177 5825 25211
rect 5859 25208 5871 25211
rect 6273 25211 6331 25217
rect 6273 25208 6285 25211
rect 5859 25180 6285 25208
rect 5859 25177 5871 25180
rect 5813 25171 5871 25177
rect 6273 25177 6285 25180
rect 6319 25177 6331 25211
rect 6273 25171 6331 25177
rect 7552 25211 7610 25217
rect 7552 25177 7564 25211
rect 7598 25208 7610 25211
rect 7742 25208 7748 25220
rect 7598 25180 7748 25208
rect 7598 25177 7610 25180
rect 7552 25171 7610 25177
rect 7742 25168 7748 25180
rect 7800 25168 7806 25220
rect 9508 25208 9536 25239
rect 8680 25180 9536 25208
rect 8570 25100 8576 25152
rect 8628 25140 8634 25152
rect 8680 25149 8708 25180
rect 8665 25143 8723 25149
rect 8665 25140 8677 25143
rect 8628 25112 8677 25140
rect 8628 25100 8634 25112
rect 8665 25109 8677 25112
rect 8711 25109 8723 25143
rect 8665 25103 8723 25109
rect 8938 25100 8944 25152
rect 8996 25100 9002 25152
rect 9306 25100 9312 25152
rect 9364 25140 9370 25152
rect 9646 25140 9674 25248
rect 9861 25245 9873 25248
rect 9907 25245 9919 25279
rect 9861 25239 9919 25245
rect 9950 25236 9956 25288
rect 10008 25236 10014 25288
rect 10244 25285 10272 25316
rect 12066 25304 12072 25356
rect 12124 25344 12130 25356
rect 12176 25344 12204 25375
rect 12805 25347 12863 25353
rect 12805 25344 12817 25347
rect 12124 25316 12817 25344
rect 12124 25304 12130 25316
rect 12805 25313 12817 25316
rect 12851 25313 12863 25347
rect 22081 25344 22109 25452
rect 22646 25440 22652 25492
rect 22704 25440 22710 25492
rect 23474 25440 23480 25492
rect 23532 25440 23538 25492
rect 23658 25440 23664 25492
rect 23716 25480 23722 25492
rect 24397 25483 24455 25489
rect 24397 25480 24409 25483
rect 23716 25452 24409 25480
rect 23716 25440 23722 25452
rect 24397 25449 24409 25452
rect 24443 25449 24455 25483
rect 24397 25443 24455 25449
rect 26050 25440 26056 25492
rect 26108 25440 26114 25492
rect 22664 25412 22692 25440
rect 22664 25384 25452 25412
rect 24026 25344 24032 25356
rect 22081 25316 24032 25344
rect 12805 25307 12863 25313
rect 24026 25304 24032 25316
rect 24084 25304 24090 25356
rect 24486 25304 24492 25356
rect 24544 25344 24550 25356
rect 25041 25347 25099 25353
rect 25041 25344 25053 25347
rect 24544 25316 25053 25344
rect 24544 25304 24550 25316
rect 25041 25313 25053 25316
rect 25087 25344 25099 25347
rect 25130 25344 25136 25356
rect 25087 25316 25136 25344
rect 25087 25313 25099 25316
rect 25041 25307 25099 25313
rect 25130 25304 25136 25316
rect 25188 25304 25194 25356
rect 10229 25279 10287 25285
rect 10229 25245 10241 25279
rect 10275 25245 10287 25279
rect 10229 25239 10287 25245
rect 10778 25236 10784 25288
rect 10836 25236 10842 25288
rect 18506 25236 18512 25288
rect 18564 25276 18570 25288
rect 19334 25276 19340 25288
rect 18564 25248 19340 25276
rect 18564 25236 18570 25248
rect 19334 25236 19340 25248
rect 19392 25276 19398 25288
rect 19429 25279 19487 25285
rect 19429 25276 19441 25279
rect 19392 25248 19441 25276
rect 19392 25236 19398 25248
rect 19429 25245 19441 25248
rect 19475 25245 19487 25279
rect 19429 25239 19487 25245
rect 19886 25236 19892 25288
rect 19944 25276 19950 25288
rect 20441 25279 20499 25285
rect 20441 25276 20453 25279
rect 19944 25248 20453 25276
rect 19944 25236 19950 25248
rect 20441 25245 20453 25248
rect 20487 25245 20499 25279
rect 20441 25239 20499 25245
rect 23845 25279 23903 25285
rect 23845 25245 23857 25279
rect 23891 25276 23903 25279
rect 24394 25276 24400 25288
rect 23891 25248 24400 25276
rect 23891 25245 23903 25248
rect 23845 25239 23903 25245
rect 24394 25236 24400 25248
rect 24452 25236 24458 25288
rect 10042 25168 10048 25220
rect 10100 25168 10106 25220
rect 11048 25211 11106 25217
rect 11048 25177 11060 25211
rect 11094 25208 11106 25211
rect 11330 25208 11336 25220
rect 11094 25180 11336 25208
rect 11094 25177 11106 25180
rect 11048 25171 11106 25177
rect 11330 25168 11336 25180
rect 11388 25168 11394 25220
rect 16482 25168 16488 25220
rect 16540 25208 16546 25220
rect 23937 25211 23995 25217
rect 23937 25208 23949 25211
rect 16540 25180 23949 25208
rect 16540 25168 16546 25180
rect 23937 25177 23949 25180
rect 23983 25177 23995 25211
rect 23937 25171 23995 25177
rect 24765 25211 24823 25217
rect 24765 25177 24777 25211
rect 24811 25208 24823 25211
rect 25317 25211 25375 25217
rect 25317 25208 25329 25211
rect 24811 25180 25329 25208
rect 24811 25177 24823 25180
rect 24765 25171 24823 25177
rect 25317 25177 25329 25180
rect 25363 25177 25375 25211
rect 25424 25208 25452 25384
rect 25774 25304 25780 25356
rect 25832 25344 25838 25356
rect 25869 25347 25927 25353
rect 25869 25344 25881 25347
rect 25832 25316 25881 25344
rect 25832 25304 25838 25316
rect 25869 25313 25881 25316
rect 25915 25313 25927 25347
rect 25869 25307 25927 25313
rect 26068 25276 26096 25440
rect 26237 25279 26295 25285
rect 26237 25276 26249 25279
rect 26068 25248 26249 25276
rect 26237 25245 26249 25248
rect 26283 25245 26295 25279
rect 26237 25239 26295 25245
rect 29730 25208 29736 25220
rect 25424 25180 29736 25208
rect 25317 25171 25375 25177
rect 9364 25112 9674 25140
rect 9364 25100 9370 25112
rect 9766 25100 9772 25152
rect 9824 25140 9830 25152
rect 10594 25140 10600 25152
rect 9824 25112 10600 25140
rect 9824 25100 9830 25112
rect 10594 25100 10600 25112
rect 10652 25100 10658 25152
rect 12250 25100 12256 25152
rect 12308 25100 12314 25152
rect 19337 25143 19395 25149
rect 19337 25109 19349 25143
rect 19383 25140 19395 25143
rect 19426 25140 19432 25152
rect 19383 25112 19432 25140
rect 19383 25109 19395 25112
rect 19337 25103 19395 25109
rect 19426 25100 19432 25112
rect 19484 25100 19490 25152
rect 20625 25143 20683 25149
rect 20625 25109 20637 25143
rect 20671 25140 20683 25143
rect 21542 25140 21548 25152
rect 20671 25112 21548 25140
rect 20671 25109 20683 25112
rect 20625 25103 20683 25109
rect 21542 25100 21548 25112
rect 21600 25100 21606 25152
rect 23952 25140 23980 25171
rect 29730 25168 29736 25180
rect 29788 25168 29794 25220
rect 24857 25143 24915 25149
rect 24857 25140 24869 25143
rect 23952 25112 24869 25140
rect 24857 25109 24869 25112
rect 24903 25140 24915 25143
rect 25498 25140 25504 25152
rect 24903 25112 25504 25140
rect 24903 25109 24915 25112
rect 24857 25103 24915 25109
rect 25498 25100 25504 25112
rect 25556 25100 25562 25152
rect 26053 25143 26111 25149
rect 26053 25109 26065 25143
rect 26099 25140 26111 25143
rect 26142 25140 26148 25152
rect 26099 25112 26148 25140
rect 26099 25109 26111 25112
rect 26053 25103 26111 25109
rect 26142 25100 26148 25112
rect 26200 25100 26206 25152
rect 1104 25050 31832 25072
rect 1104 24998 4922 25050
rect 4974 24998 4986 25050
rect 5038 24998 5050 25050
rect 5102 24998 5114 25050
rect 5166 24998 5178 25050
rect 5230 24998 5242 25050
rect 5294 24998 10922 25050
rect 10974 24998 10986 25050
rect 11038 24998 11050 25050
rect 11102 24998 11114 25050
rect 11166 24998 11178 25050
rect 11230 24998 11242 25050
rect 11294 24998 16922 25050
rect 16974 24998 16986 25050
rect 17038 24998 17050 25050
rect 17102 24998 17114 25050
rect 17166 24998 17178 25050
rect 17230 24998 17242 25050
rect 17294 24998 22922 25050
rect 22974 24998 22986 25050
rect 23038 24998 23050 25050
rect 23102 24998 23114 25050
rect 23166 24998 23178 25050
rect 23230 24998 23242 25050
rect 23294 24998 28922 25050
rect 28974 24998 28986 25050
rect 29038 24998 29050 25050
rect 29102 24998 29114 25050
rect 29166 24998 29178 25050
rect 29230 24998 29242 25050
rect 29294 24998 31832 25050
rect 1104 24976 31832 24998
rect 4798 24896 4804 24948
rect 4856 24936 4862 24948
rect 5353 24939 5411 24945
rect 5353 24936 5365 24939
rect 4856 24908 5365 24936
rect 4856 24896 4862 24908
rect 5353 24905 5365 24908
rect 5399 24905 5411 24939
rect 5353 24899 5411 24905
rect 5534 24896 5540 24948
rect 5592 24896 5598 24948
rect 7742 24896 7748 24948
rect 7800 24896 7806 24948
rect 8389 24939 8447 24945
rect 8389 24905 8401 24939
rect 8435 24936 8447 24939
rect 8938 24936 8944 24948
rect 8435 24908 8944 24936
rect 8435 24905 8447 24908
rect 8389 24899 8447 24905
rect 8938 24896 8944 24908
rect 8996 24896 9002 24948
rect 11149 24939 11207 24945
rect 11149 24905 11161 24939
rect 11195 24936 11207 24939
rect 11330 24936 11336 24948
rect 11195 24908 11336 24936
rect 11195 24905 11207 24908
rect 11149 24899 11207 24905
rect 11330 24896 11336 24908
rect 11388 24896 11394 24948
rect 11885 24939 11943 24945
rect 11885 24905 11897 24939
rect 11931 24936 11943 24939
rect 12250 24936 12256 24948
rect 11931 24908 12256 24936
rect 11931 24905 11943 24908
rect 11885 24899 11943 24905
rect 12250 24896 12256 24908
rect 12308 24896 12314 24948
rect 16482 24936 16488 24948
rect 13464 24908 16488 24936
rect 4148 24871 4206 24877
rect 4148 24837 4160 24871
rect 4194 24868 4206 24871
rect 4614 24868 4620 24880
rect 4194 24840 4620 24868
rect 4194 24837 4206 24840
rect 4148 24831 4206 24837
rect 4614 24828 4620 24840
rect 4672 24828 4678 24880
rect 3881 24803 3939 24809
rect 3881 24769 3893 24803
rect 3927 24800 3939 24803
rect 3970 24800 3976 24812
rect 3927 24772 3976 24800
rect 3927 24769 3939 24772
rect 3881 24763 3939 24769
rect 3970 24760 3976 24772
rect 4028 24760 4034 24812
rect 5552 24809 5580 24896
rect 5537 24803 5595 24809
rect 5537 24769 5549 24803
rect 5583 24769 5595 24803
rect 5537 24763 5595 24769
rect 7929 24803 7987 24809
rect 7929 24769 7941 24803
rect 7975 24800 7987 24803
rect 8846 24800 8852 24812
rect 7975 24772 8064 24800
rect 7975 24769 7987 24772
rect 7929 24763 7987 24769
rect 934 24692 940 24744
rect 992 24732 998 24744
rect 1397 24735 1455 24741
rect 1397 24732 1409 24735
rect 992 24704 1409 24732
rect 992 24692 998 24704
rect 1397 24701 1409 24704
rect 1443 24701 1455 24735
rect 1397 24695 1455 24701
rect 1673 24735 1731 24741
rect 1673 24701 1685 24735
rect 1719 24732 1731 24735
rect 3786 24732 3792 24744
rect 1719 24704 3792 24732
rect 1719 24701 1731 24704
rect 1673 24695 1731 24701
rect 3786 24692 3792 24704
rect 3844 24692 3850 24744
rect 5261 24667 5319 24673
rect 5261 24633 5273 24667
rect 5307 24664 5319 24667
rect 6914 24664 6920 24676
rect 5307 24636 6920 24664
rect 5307 24633 5319 24636
rect 5261 24627 5319 24633
rect 6914 24624 6920 24636
rect 6972 24624 6978 24676
rect 8036 24673 8064 24772
rect 8588 24772 8852 24800
rect 8294 24692 8300 24744
rect 8352 24732 8358 24744
rect 8588 24741 8616 24772
rect 8846 24760 8852 24772
rect 8904 24760 8910 24812
rect 10873 24803 10931 24809
rect 10873 24800 10885 24803
rect 10350 24772 10885 24800
rect 10873 24769 10885 24772
rect 10919 24769 10931 24803
rect 10873 24763 10931 24769
rect 10965 24803 11023 24809
rect 10965 24769 10977 24803
rect 11011 24769 11023 24803
rect 10965 24763 11023 24769
rect 11333 24803 11391 24809
rect 11333 24769 11345 24803
rect 11379 24800 11391 24803
rect 11977 24803 12035 24809
rect 11379 24772 11560 24800
rect 11379 24769 11391 24772
rect 11333 24763 11391 24769
rect 8481 24735 8539 24741
rect 8481 24732 8493 24735
rect 8352 24704 8493 24732
rect 8352 24692 8358 24704
rect 8481 24701 8493 24704
rect 8527 24701 8539 24735
rect 8481 24695 8539 24701
rect 8573 24735 8631 24741
rect 8573 24701 8585 24735
rect 8619 24701 8631 24735
rect 8573 24695 8631 24701
rect 8021 24667 8079 24673
rect 8021 24633 8033 24667
rect 8067 24633 8079 24667
rect 8496 24664 8524 24695
rect 8662 24692 8668 24744
rect 8720 24732 8726 24744
rect 8941 24735 8999 24741
rect 8941 24732 8953 24735
rect 8720 24704 8953 24732
rect 8720 24692 8726 24704
rect 8941 24701 8953 24704
rect 8987 24701 8999 24735
rect 8941 24695 8999 24701
rect 9214 24692 9220 24744
rect 9272 24692 9278 24744
rect 10980 24732 11008 24763
rect 10612 24704 11008 24732
rect 10612 24676 10640 24704
rect 8496 24636 8616 24664
rect 8021 24627 8079 24633
rect 8588 24596 8616 24636
rect 10594 24624 10600 24676
rect 10652 24624 10658 24676
rect 10686 24624 10692 24676
rect 10744 24624 10750 24676
rect 11532 24673 11560 24772
rect 11977 24769 11989 24803
rect 12023 24800 12035 24803
rect 13464 24800 13492 24908
rect 16482 24896 16488 24908
rect 16540 24896 16546 24948
rect 19886 24896 19892 24948
rect 19944 24896 19950 24948
rect 25774 24936 25780 24948
rect 25424 24908 25780 24936
rect 19426 24828 19432 24880
rect 19484 24828 19490 24880
rect 24302 24828 24308 24880
rect 24360 24868 24366 24880
rect 24489 24871 24547 24877
rect 24489 24868 24501 24871
rect 24360 24840 24501 24868
rect 24360 24828 24366 24840
rect 24489 24837 24501 24840
rect 24535 24837 24547 24871
rect 24489 24831 24547 24837
rect 12023 24772 13492 24800
rect 14001 24803 14059 24809
rect 12023 24769 12035 24772
rect 11977 24763 12035 24769
rect 14001 24769 14013 24803
rect 14047 24800 14059 24803
rect 14826 24800 14832 24812
rect 14047 24772 14832 24800
rect 14047 24769 14059 24772
rect 14001 24763 14059 24769
rect 11517 24667 11575 24673
rect 11517 24633 11529 24667
rect 11563 24633 11575 24667
rect 11517 24627 11575 24633
rect 9674 24596 9680 24608
rect 8588 24568 9680 24596
rect 9674 24556 9680 24568
rect 9732 24596 9738 24608
rect 11992 24596 12020 24763
rect 14826 24760 14832 24772
rect 14884 24760 14890 24812
rect 20070 24760 20076 24812
rect 20128 24760 20134 24812
rect 24210 24760 24216 24812
rect 24268 24760 24274 24812
rect 25424 24809 25452 24908
rect 25774 24896 25780 24908
rect 25832 24896 25838 24948
rect 29362 24896 29368 24948
rect 29420 24936 29426 24948
rect 29641 24939 29699 24945
rect 29641 24936 29653 24939
rect 29420 24908 29653 24936
rect 29420 24896 29426 24908
rect 29641 24905 29653 24908
rect 29687 24905 29699 24939
rect 29641 24899 29699 24905
rect 28810 24828 28816 24880
rect 28868 24868 28874 24880
rect 29454 24868 29460 24880
rect 28868 24840 29460 24868
rect 28868 24828 28874 24840
rect 29454 24828 29460 24840
rect 29512 24828 29518 24880
rect 29549 24871 29607 24877
rect 29549 24837 29561 24871
rect 29595 24868 29607 24871
rect 30285 24871 30343 24877
rect 30285 24868 30297 24871
rect 29595 24840 30297 24868
rect 29595 24837 29607 24840
rect 29549 24831 29607 24837
rect 30285 24837 30297 24840
rect 30331 24837 30343 24871
rect 30285 24831 30343 24837
rect 24397 24803 24455 24809
rect 24397 24769 24409 24803
rect 24443 24769 24455 24803
rect 24397 24763 24455 24769
rect 24581 24803 24639 24809
rect 24581 24769 24593 24803
rect 24627 24769 24639 24803
rect 24581 24763 24639 24769
rect 25409 24803 25467 24809
rect 25409 24769 25421 24803
rect 25455 24769 25467 24803
rect 25409 24763 25467 24769
rect 25593 24803 25651 24809
rect 25593 24769 25605 24803
rect 25639 24769 25651 24803
rect 25593 24763 25651 24769
rect 25685 24803 25743 24809
rect 25685 24769 25697 24803
rect 25731 24769 25743 24803
rect 25685 24763 25743 24769
rect 25777 24803 25835 24809
rect 25777 24769 25789 24803
rect 25823 24800 25835 24803
rect 26510 24800 26516 24812
rect 25823 24772 26516 24800
rect 25823 24769 25835 24772
rect 25777 24763 25835 24769
rect 12158 24692 12164 24744
rect 12216 24692 12222 24744
rect 13725 24735 13783 24741
rect 13725 24701 13737 24735
rect 13771 24732 13783 24735
rect 13814 24732 13820 24744
rect 13771 24704 13820 24732
rect 13771 24701 13783 24704
rect 13725 24695 13783 24701
rect 13814 24692 13820 24704
rect 13872 24692 13878 24744
rect 17954 24692 17960 24744
rect 18012 24732 18018 24744
rect 18141 24735 18199 24741
rect 18141 24732 18153 24735
rect 18012 24704 18153 24732
rect 18012 24692 18018 24704
rect 18141 24701 18153 24704
rect 18187 24701 18199 24735
rect 18141 24695 18199 24701
rect 18414 24692 18420 24744
rect 18472 24692 18478 24744
rect 24118 24692 24124 24744
rect 24176 24732 24182 24744
rect 24412 24732 24440 24763
rect 24176 24704 24440 24732
rect 24176 24692 24182 24704
rect 13909 24667 13967 24673
rect 13909 24633 13921 24667
rect 13955 24664 13967 24667
rect 13998 24664 14004 24676
rect 13955 24636 14004 24664
rect 13955 24633 13967 24636
rect 13909 24627 13967 24633
rect 13998 24624 14004 24636
rect 14056 24624 14062 24676
rect 24302 24624 24308 24676
rect 24360 24664 24366 24676
rect 24596 24664 24624 24763
rect 24360 24636 24624 24664
rect 25608 24664 25636 24763
rect 25700 24732 25728 24763
rect 26510 24760 26516 24772
rect 26568 24760 26574 24812
rect 27154 24760 27160 24812
rect 27212 24760 27218 24812
rect 27246 24760 27252 24812
rect 27304 24760 27310 24812
rect 27338 24760 27344 24812
rect 27396 24760 27402 24812
rect 27522 24760 27528 24812
rect 27580 24760 27586 24812
rect 29362 24760 29368 24812
rect 29420 24800 29426 24812
rect 30009 24803 30067 24809
rect 30009 24800 30021 24803
rect 29420 24772 30021 24800
rect 29420 24760 29426 24772
rect 30009 24769 30021 24772
rect 30055 24769 30067 24803
rect 30009 24763 30067 24769
rect 26878 24732 26884 24744
rect 25700 24704 26884 24732
rect 26878 24692 26884 24704
rect 26936 24692 26942 24744
rect 28537 24735 28595 24741
rect 28537 24701 28549 24735
rect 28583 24732 28595 24735
rect 28718 24732 28724 24744
rect 28583 24704 28724 24732
rect 28583 24701 28595 24704
rect 28537 24695 28595 24701
rect 28718 24692 28724 24704
rect 28776 24692 28782 24744
rect 29730 24692 29736 24744
rect 29788 24692 29794 24744
rect 30837 24735 30895 24741
rect 30837 24701 30849 24735
rect 30883 24701 30895 24735
rect 30837 24695 30895 24701
rect 26694 24664 26700 24676
rect 25608 24636 26700 24664
rect 24360 24624 24366 24636
rect 26694 24624 26700 24636
rect 26752 24624 26758 24676
rect 30852 24608 30880 24695
rect 9732 24568 12020 24596
rect 9732 24556 9738 24568
rect 12158 24556 12164 24608
rect 12216 24596 12222 24608
rect 13817 24599 13875 24605
rect 13817 24596 13829 24599
rect 12216 24568 13829 24596
rect 12216 24556 12222 24568
rect 13817 24565 13829 24568
rect 13863 24596 13875 24599
rect 14090 24596 14096 24608
rect 13863 24568 14096 24596
rect 13863 24565 13875 24568
rect 13817 24559 13875 24565
rect 14090 24556 14096 24568
rect 14148 24556 14154 24608
rect 19426 24556 19432 24608
rect 19484 24596 19490 24608
rect 20165 24599 20223 24605
rect 20165 24596 20177 24599
rect 19484 24568 20177 24596
rect 19484 24556 19490 24568
rect 20165 24565 20177 24568
rect 20211 24565 20223 24599
rect 20165 24559 20223 24565
rect 24762 24556 24768 24608
rect 24820 24556 24826 24608
rect 25958 24556 25964 24608
rect 26016 24556 26022 24608
rect 26970 24556 26976 24608
rect 27028 24556 27034 24608
rect 28994 24556 29000 24608
rect 29052 24596 29058 24608
rect 29089 24599 29147 24605
rect 29089 24596 29101 24599
rect 29052 24568 29101 24596
rect 29052 24556 29058 24568
rect 29089 24565 29101 24568
rect 29135 24565 29147 24599
rect 29089 24559 29147 24565
rect 29178 24556 29184 24608
rect 29236 24556 29242 24608
rect 30190 24556 30196 24608
rect 30248 24556 30254 24608
rect 30834 24556 30840 24608
rect 30892 24556 30898 24608
rect 1104 24506 31832 24528
rect 1104 24454 4182 24506
rect 4234 24454 4246 24506
rect 4298 24454 4310 24506
rect 4362 24454 4374 24506
rect 4426 24454 4438 24506
rect 4490 24454 4502 24506
rect 4554 24454 10182 24506
rect 10234 24454 10246 24506
rect 10298 24454 10310 24506
rect 10362 24454 10374 24506
rect 10426 24454 10438 24506
rect 10490 24454 10502 24506
rect 10554 24454 16182 24506
rect 16234 24454 16246 24506
rect 16298 24454 16310 24506
rect 16362 24454 16374 24506
rect 16426 24454 16438 24506
rect 16490 24454 16502 24506
rect 16554 24454 22182 24506
rect 22234 24454 22246 24506
rect 22298 24454 22310 24506
rect 22362 24454 22374 24506
rect 22426 24454 22438 24506
rect 22490 24454 22502 24506
rect 22554 24454 28182 24506
rect 28234 24454 28246 24506
rect 28298 24454 28310 24506
rect 28362 24454 28374 24506
rect 28426 24454 28438 24506
rect 28490 24454 28502 24506
rect 28554 24454 31832 24506
rect 1104 24432 31832 24454
rect 9214 24352 9220 24404
rect 9272 24392 9278 24404
rect 9309 24395 9367 24401
rect 9309 24392 9321 24395
rect 9272 24364 9321 24392
rect 9272 24352 9278 24364
rect 9309 24361 9321 24364
rect 9355 24361 9367 24395
rect 9309 24355 9367 24361
rect 9490 24352 9496 24404
rect 9548 24392 9554 24404
rect 12158 24392 12164 24404
rect 9548 24364 12164 24392
rect 9548 24352 9554 24364
rect 12158 24352 12164 24364
rect 12216 24352 12222 24404
rect 12342 24352 12348 24404
rect 12400 24392 12406 24404
rect 15654 24392 15660 24404
rect 12400 24364 15660 24392
rect 12400 24352 12406 24364
rect 15654 24352 15660 24364
rect 15712 24352 15718 24404
rect 16669 24395 16727 24401
rect 16669 24361 16681 24395
rect 16715 24392 16727 24395
rect 18414 24392 18420 24404
rect 16715 24364 18420 24392
rect 16715 24361 16727 24364
rect 16669 24355 16727 24361
rect 18414 24352 18420 24364
rect 18472 24352 18478 24404
rect 18874 24352 18880 24404
rect 18932 24352 18938 24404
rect 20070 24352 20076 24404
rect 20128 24352 20134 24404
rect 21560 24364 21772 24392
rect 6089 24327 6147 24333
rect 6089 24293 6101 24327
rect 6135 24324 6147 24327
rect 8481 24327 8539 24333
rect 6135 24296 6914 24324
rect 6135 24293 6147 24296
rect 6089 24287 6147 24293
rect 6886 24256 6914 24296
rect 8481 24293 8493 24327
rect 8527 24324 8539 24327
rect 11425 24327 11483 24333
rect 11425 24324 11437 24327
rect 8527 24296 11437 24324
rect 8527 24293 8539 24296
rect 8481 24287 8539 24293
rect 11425 24293 11437 24296
rect 11471 24293 11483 24327
rect 21560 24324 21588 24364
rect 11425 24287 11483 24293
rect 12406 24296 21588 24324
rect 21744 24324 21772 24364
rect 25958 24352 25964 24404
rect 26016 24352 26022 24404
rect 26970 24352 26976 24404
rect 27028 24352 27034 24404
rect 29178 24352 29184 24404
rect 29236 24352 29242 24404
rect 29362 24352 29368 24404
rect 29420 24352 29426 24404
rect 26237 24327 26295 24333
rect 26237 24324 26249 24327
rect 21744 24296 26249 24324
rect 10321 24259 10379 24265
rect 6886 24228 8340 24256
rect 5537 24191 5595 24197
rect 5537 24157 5549 24191
rect 5583 24188 5595 24191
rect 5626 24188 5632 24200
rect 5583 24160 5632 24188
rect 5583 24157 5595 24160
rect 5537 24151 5595 24157
rect 5626 24148 5632 24160
rect 5684 24148 5690 24200
rect 5902 24148 5908 24200
rect 5960 24148 5966 24200
rect 8312 24197 8340 24228
rect 10321 24225 10333 24259
rect 10367 24256 10379 24259
rect 11793 24259 11851 24265
rect 11793 24256 11805 24259
rect 10367 24228 10824 24256
rect 10367 24225 10379 24228
rect 10321 24219 10379 24225
rect 8021 24191 8079 24197
rect 8021 24157 8033 24191
rect 8067 24157 8079 24191
rect 8021 24151 8079 24157
rect 8297 24191 8355 24197
rect 8297 24157 8309 24191
rect 8343 24157 8355 24191
rect 8297 24151 8355 24157
rect 9493 24191 9551 24197
rect 9493 24157 9505 24191
rect 9539 24188 9551 24191
rect 10045 24191 10103 24197
rect 9539 24160 9720 24188
rect 9539 24157 9551 24160
rect 9493 24151 9551 24157
rect 5718 24080 5724 24132
rect 5776 24080 5782 24132
rect 5813 24123 5871 24129
rect 5813 24089 5825 24123
rect 5859 24120 5871 24123
rect 6914 24120 6920 24132
rect 5859 24092 6920 24120
rect 5859 24089 5871 24092
rect 5813 24083 5871 24089
rect 6914 24080 6920 24092
rect 6972 24080 6978 24132
rect 8036 24064 8064 24151
rect 8113 24123 8171 24129
rect 8113 24089 8125 24123
rect 8159 24120 8171 24123
rect 8570 24120 8576 24132
rect 8159 24092 8576 24120
rect 8159 24089 8171 24092
rect 8113 24083 8171 24089
rect 8570 24080 8576 24092
rect 8628 24080 8634 24132
rect 8018 24012 8024 24064
rect 8076 24012 8082 24064
rect 9692 24061 9720 24160
rect 10045 24157 10057 24191
rect 10091 24188 10103 24191
rect 10686 24188 10692 24200
rect 10091 24160 10692 24188
rect 10091 24157 10103 24160
rect 10045 24151 10103 24157
rect 10686 24148 10692 24160
rect 10744 24148 10750 24200
rect 10796 24120 10824 24228
rect 11256 24228 11805 24256
rect 11256 24197 11284 24228
rect 11793 24225 11805 24228
rect 11839 24225 11851 24259
rect 11793 24219 11851 24225
rect 11241 24191 11299 24197
rect 11241 24157 11253 24191
rect 11287 24157 11299 24191
rect 11241 24151 11299 24157
rect 11333 24191 11391 24197
rect 11333 24157 11345 24191
rect 11379 24188 11391 24191
rect 11422 24188 11428 24200
rect 11379 24160 11428 24188
rect 11379 24157 11391 24160
rect 11333 24151 11391 24157
rect 11422 24148 11428 24160
rect 11480 24148 11486 24200
rect 11517 24191 11575 24197
rect 11517 24157 11529 24191
rect 11563 24188 11575 24191
rect 12406 24188 12434 24296
rect 26237 24293 26249 24296
rect 26283 24293 26295 24327
rect 26237 24287 26295 24293
rect 13998 24256 14004 24268
rect 13464 24228 14004 24256
rect 11563 24160 12434 24188
rect 11563 24157 11575 24160
rect 11517 24151 11575 24157
rect 12986 24148 12992 24200
rect 13044 24188 13050 24200
rect 13464 24197 13492 24228
rect 13998 24216 14004 24228
rect 14056 24256 14062 24268
rect 14056 24228 14780 24256
rect 14056 24216 14062 24228
rect 14752 24200 14780 24228
rect 16298 24216 16304 24268
rect 16356 24216 16362 24268
rect 19610 24216 19616 24268
rect 19668 24256 19674 24268
rect 19914 24259 19972 24265
rect 19914 24256 19926 24259
rect 19668 24228 19926 24256
rect 19668 24216 19674 24228
rect 19914 24225 19926 24228
rect 19960 24256 19972 24259
rect 20530 24256 20536 24268
rect 19960 24228 20536 24256
rect 19960 24225 19972 24228
rect 19914 24219 19972 24225
rect 20530 24216 20536 24228
rect 20588 24256 20594 24268
rect 21174 24256 21180 24268
rect 20588 24228 21180 24256
rect 20588 24216 20594 24228
rect 21174 24216 21180 24228
rect 21232 24256 21238 24268
rect 21361 24259 21419 24265
rect 21361 24256 21373 24259
rect 21232 24228 21373 24256
rect 21232 24216 21238 24228
rect 21361 24225 21373 24228
rect 21407 24225 21419 24259
rect 21361 24219 21419 24225
rect 24762 24216 24768 24268
rect 24820 24216 24826 24268
rect 25961 24259 26019 24265
rect 25961 24225 25973 24259
rect 26007 24256 26019 24259
rect 26988 24256 27016 24352
rect 29196 24324 29224 24352
rect 26007 24228 27016 24256
rect 28368 24296 29224 24324
rect 26007 24225 26019 24228
rect 25961 24219 26019 24225
rect 13449 24191 13507 24197
rect 13449 24188 13461 24191
rect 13044 24160 13461 24188
rect 13044 24148 13050 24160
rect 13449 24157 13461 24160
rect 13495 24157 13507 24191
rect 13449 24151 13507 24157
rect 14090 24148 14096 24200
rect 14148 24188 14154 24200
rect 14645 24191 14703 24197
rect 14645 24188 14657 24191
rect 14148 24160 14657 24188
rect 14148 24148 14154 24160
rect 14645 24157 14657 24160
rect 14691 24157 14703 24191
rect 14645 24151 14703 24157
rect 14734 24148 14740 24200
rect 14792 24188 14798 24200
rect 15013 24191 15071 24197
rect 15013 24188 15025 24191
rect 14792 24160 15025 24188
rect 14792 24148 14798 24160
rect 15013 24157 15025 24160
rect 15059 24188 15071 24191
rect 16393 24191 16451 24197
rect 16393 24188 16405 24191
rect 15059 24160 16405 24188
rect 15059 24157 15071 24160
rect 15013 24151 15071 24157
rect 16393 24157 16405 24160
rect 16439 24157 16451 24191
rect 16393 24151 16451 24157
rect 18969 24191 19027 24197
rect 18969 24157 18981 24191
rect 19015 24188 19027 24191
rect 19058 24188 19064 24200
rect 19015 24160 19064 24188
rect 19015 24157 19027 24160
rect 18969 24151 19027 24157
rect 10704 24092 10824 24120
rect 11977 24123 12035 24129
rect 10704 24064 10732 24092
rect 11977 24089 11989 24123
rect 12023 24120 12035 24123
rect 12066 24120 12072 24132
rect 12023 24092 12072 24120
rect 12023 24089 12035 24092
rect 11977 24083 12035 24089
rect 12066 24080 12072 24092
rect 12124 24080 12130 24132
rect 12158 24080 12164 24132
rect 12216 24080 12222 24132
rect 13265 24123 13323 24129
rect 13265 24089 13277 24123
rect 13311 24120 13323 24123
rect 13817 24123 13875 24129
rect 13311 24092 13768 24120
rect 13311 24089 13323 24092
rect 13265 24083 13323 24089
rect 9677 24055 9735 24061
rect 9677 24021 9689 24055
rect 9723 24021 9735 24055
rect 9677 24015 9735 24021
rect 9950 24012 9956 24064
rect 10008 24052 10014 24064
rect 10137 24055 10195 24061
rect 10137 24052 10149 24055
rect 10008 24024 10149 24052
rect 10008 24012 10014 24024
rect 10137 24021 10149 24024
rect 10183 24021 10195 24055
rect 10137 24015 10195 24021
rect 10686 24012 10692 24064
rect 10744 24012 10750 24064
rect 11701 24055 11759 24061
rect 11701 24021 11713 24055
rect 11747 24052 11759 24055
rect 12710 24052 12716 24064
rect 11747 24024 12716 24052
rect 11747 24021 11759 24024
rect 11701 24015 11759 24021
rect 12710 24012 12716 24024
rect 12768 24012 12774 24064
rect 13538 24012 13544 24064
rect 13596 24012 13602 24064
rect 13630 24012 13636 24064
rect 13688 24012 13694 24064
rect 13740 24052 13768 24092
rect 13817 24089 13829 24123
rect 13863 24120 13875 24123
rect 14185 24123 14243 24129
rect 14185 24120 14197 24123
rect 13863 24092 14197 24120
rect 13863 24089 13875 24092
rect 13817 24083 13875 24089
rect 14185 24089 14197 24092
rect 14231 24089 14243 24123
rect 16408 24120 16436 24151
rect 19058 24148 19064 24160
rect 19116 24148 19122 24200
rect 19429 24191 19487 24197
rect 19429 24157 19441 24191
rect 19475 24188 19487 24191
rect 19518 24188 19524 24200
rect 19475 24160 19524 24188
rect 19475 24157 19487 24160
rect 19429 24151 19487 24157
rect 19518 24148 19524 24160
rect 19576 24188 19582 24200
rect 20070 24188 20076 24200
rect 19576 24160 20076 24188
rect 19576 24148 19582 24160
rect 20070 24148 20076 24160
rect 20128 24188 20134 24200
rect 20257 24191 20315 24197
rect 20257 24188 20269 24191
rect 20128 24160 20269 24188
rect 20128 24148 20134 24160
rect 20257 24157 20269 24160
rect 20303 24157 20315 24191
rect 20257 24151 20315 24157
rect 20346 24148 20352 24200
rect 20404 24148 20410 24200
rect 20438 24148 20444 24200
rect 20496 24148 20502 24200
rect 21450 24148 21456 24200
rect 21508 24148 21514 24200
rect 21542 24148 21548 24200
rect 21600 24148 21606 24200
rect 21637 24191 21695 24197
rect 21637 24157 21649 24191
rect 21683 24157 21695 24191
rect 21637 24151 21695 24157
rect 22925 24191 22983 24197
rect 22925 24157 22937 24191
rect 22971 24157 22983 24191
rect 22925 24151 22983 24157
rect 23201 24191 23259 24197
rect 23201 24157 23213 24191
rect 23247 24188 23259 24191
rect 23382 24188 23388 24200
rect 23247 24160 23388 24188
rect 23247 24157 23259 24160
rect 23201 24151 23259 24157
rect 20364 24120 20392 24148
rect 16408 24092 20392 24120
rect 14185 24083 14243 24089
rect 13906 24052 13912 24064
rect 13740 24024 13912 24052
rect 13906 24012 13912 24024
rect 13964 24012 13970 24064
rect 14274 24012 14280 24064
rect 14332 24012 14338 24064
rect 14458 24012 14464 24064
rect 14516 24052 14522 24064
rect 14829 24055 14887 24061
rect 14829 24052 14841 24055
rect 14516 24024 14841 24052
rect 14516 24012 14522 24024
rect 14829 24021 14841 24024
rect 14875 24021 14887 24055
rect 14829 24015 14887 24021
rect 15105 24055 15163 24061
rect 15105 24021 15117 24055
rect 15151 24052 15163 24055
rect 15286 24052 15292 24064
rect 15151 24024 15292 24052
rect 15151 24021 15163 24024
rect 15105 24015 15163 24021
rect 15286 24012 15292 24024
rect 15344 24012 15350 24064
rect 19702 24012 19708 24064
rect 19760 24012 19766 24064
rect 19797 24055 19855 24061
rect 19797 24021 19809 24055
rect 19843 24052 19855 24055
rect 19978 24052 19984 24064
rect 19843 24024 19984 24052
rect 19843 24021 19855 24024
rect 19797 24015 19855 24021
rect 19978 24012 19984 24024
rect 20036 24052 20042 24064
rect 20456 24052 20484 24148
rect 20714 24080 20720 24132
rect 20772 24080 20778 24132
rect 21652 24120 21680 24151
rect 21560 24092 21680 24120
rect 21821 24123 21879 24129
rect 21560 24052 21588 24092
rect 21821 24089 21833 24123
rect 21867 24120 21879 24123
rect 22940 24120 22968 24151
rect 23382 24148 23388 24160
rect 23440 24148 23446 24200
rect 24780 24188 24808 24216
rect 25777 24191 25835 24197
rect 25777 24188 25789 24191
rect 24780 24160 25789 24188
rect 25777 24157 25789 24160
rect 25823 24157 25835 24191
rect 25777 24151 25835 24157
rect 26050 24148 26056 24200
rect 26108 24148 26114 24200
rect 28368 24197 28396 24296
rect 28810 24216 28816 24268
rect 28868 24216 28874 24268
rect 28905 24259 28963 24265
rect 28905 24225 28917 24259
rect 28951 24256 28963 24259
rect 29270 24256 29276 24268
rect 28951 24228 29276 24256
rect 28951 24225 28963 24228
rect 28905 24219 28963 24225
rect 29270 24216 29276 24228
rect 29328 24216 29334 24268
rect 28353 24191 28411 24197
rect 28353 24157 28365 24191
rect 28399 24157 28411 24191
rect 29549 24191 29607 24197
rect 29549 24188 29561 24191
rect 28353 24151 28411 24157
rect 28828 24160 29561 24188
rect 28828 24132 28856 24160
rect 29549 24157 29561 24160
rect 29595 24157 29607 24191
rect 29549 24151 29607 24157
rect 24949 24123 25007 24129
rect 24949 24120 24961 24123
rect 21867 24092 24961 24120
rect 21867 24089 21879 24092
rect 21821 24083 21879 24089
rect 24949 24089 24961 24092
rect 24995 24089 25007 24123
rect 24949 24083 25007 24089
rect 25133 24123 25191 24129
rect 25133 24089 25145 24123
rect 25179 24089 25191 24123
rect 25133 24083 25191 24089
rect 20036 24024 21588 24052
rect 25148 24052 25176 24083
rect 28810 24080 28816 24132
rect 28868 24080 28874 24132
rect 28994 24080 29000 24132
rect 29052 24080 29058 24132
rect 29794 24123 29852 24129
rect 29794 24120 29806 24123
rect 29196 24092 29806 24120
rect 26510 24052 26516 24064
rect 25148 24024 26516 24052
rect 20036 24012 20042 24024
rect 26510 24012 26516 24024
rect 26568 24012 26574 24064
rect 28537 24055 28595 24061
rect 28537 24021 28549 24055
rect 28583 24052 28595 24055
rect 29196 24052 29224 24092
rect 29794 24089 29806 24092
rect 29840 24089 29852 24123
rect 29794 24083 29852 24089
rect 28583 24024 29224 24052
rect 28583 24021 28595 24024
rect 28537 24015 28595 24021
rect 29546 24012 29552 24064
rect 29604 24052 29610 24064
rect 30834 24052 30840 24064
rect 29604 24024 30840 24052
rect 29604 24012 29610 24024
rect 30834 24012 30840 24024
rect 30892 24052 30898 24064
rect 30929 24055 30987 24061
rect 30929 24052 30941 24055
rect 30892 24024 30941 24052
rect 30892 24012 30898 24024
rect 30929 24021 30941 24024
rect 30975 24021 30987 24055
rect 30929 24015 30987 24021
rect 1104 23962 31832 23984
rect 1104 23910 4922 23962
rect 4974 23910 4986 23962
rect 5038 23910 5050 23962
rect 5102 23910 5114 23962
rect 5166 23910 5178 23962
rect 5230 23910 5242 23962
rect 5294 23910 10922 23962
rect 10974 23910 10986 23962
rect 11038 23910 11050 23962
rect 11102 23910 11114 23962
rect 11166 23910 11178 23962
rect 11230 23910 11242 23962
rect 11294 23910 16922 23962
rect 16974 23910 16986 23962
rect 17038 23910 17050 23962
rect 17102 23910 17114 23962
rect 17166 23910 17178 23962
rect 17230 23910 17242 23962
rect 17294 23910 22922 23962
rect 22974 23910 22986 23962
rect 23038 23910 23050 23962
rect 23102 23910 23114 23962
rect 23166 23910 23178 23962
rect 23230 23910 23242 23962
rect 23294 23910 28922 23962
rect 28974 23910 28986 23962
rect 29038 23910 29050 23962
rect 29102 23910 29114 23962
rect 29166 23910 29178 23962
rect 29230 23910 29242 23962
rect 29294 23910 31832 23962
rect 1104 23888 31832 23910
rect 3786 23808 3792 23860
rect 3844 23848 3850 23860
rect 12526 23848 12532 23860
rect 3844 23820 12532 23848
rect 3844 23808 3850 23820
rect 12526 23808 12532 23820
rect 12584 23808 12590 23860
rect 13446 23808 13452 23860
rect 13504 23848 13510 23860
rect 13504 23820 13768 23848
rect 13504 23808 13510 23820
rect 9766 23740 9772 23792
rect 9824 23780 9830 23792
rect 10042 23780 10048 23792
rect 9824 23752 10048 23780
rect 9824 23740 9830 23752
rect 10042 23740 10048 23752
rect 10100 23780 10106 23792
rect 13740 23789 13768 23820
rect 14366 23808 14372 23860
rect 14424 23848 14430 23860
rect 15933 23851 15991 23857
rect 14424 23820 14596 23848
rect 14424 23808 14430 23820
rect 14568 23789 14596 23820
rect 15120 23820 15608 23848
rect 13633 23783 13691 23789
rect 13633 23780 13645 23783
rect 10100 23752 13645 23780
rect 10100 23740 10106 23752
rect 13633 23749 13645 23752
rect 13679 23749 13691 23783
rect 13633 23743 13691 23749
rect 13725 23783 13783 23789
rect 13725 23749 13737 23783
rect 13771 23749 13783 23783
rect 13725 23743 13783 23749
rect 14553 23783 14611 23789
rect 14553 23749 14565 23783
rect 14599 23749 14611 23783
rect 14553 23743 14611 23749
rect 14642 23740 14648 23792
rect 14700 23780 14706 23792
rect 14826 23780 14832 23792
rect 14700 23752 14832 23780
rect 14700 23740 14706 23752
rect 14826 23740 14832 23752
rect 14884 23780 14890 23792
rect 15120 23780 15148 23820
rect 15580 23789 15608 23820
rect 15933 23817 15945 23851
rect 15979 23848 15991 23851
rect 16022 23848 16028 23860
rect 15979 23820 16028 23848
rect 15979 23817 15991 23820
rect 15933 23811 15991 23817
rect 16022 23808 16028 23820
rect 16080 23848 16086 23860
rect 16298 23848 16304 23860
rect 16080 23820 16304 23848
rect 16080 23808 16086 23820
rect 16298 23808 16304 23820
rect 16356 23808 16362 23860
rect 19245 23851 19303 23857
rect 19245 23817 19257 23851
rect 19291 23848 19303 23851
rect 20346 23848 20352 23860
rect 19291 23820 20352 23848
rect 19291 23817 19303 23820
rect 19245 23811 19303 23817
rect 20346 23808 20352 23820
rect 20404 23808 20410 23860
rect 20714 23808 20720 23860
rect 20772 23808 20778 23860
rect 20990 23808 20996 23860
rect 21048 23848 21054 23860
rect 24302 23848 24308 23860
rect 21048 23820 24308 23848
rect 21048 23808 21054 23820
rect 24302 23808 24308 23820
rect 24360 23808 24366 23860
rect 26050 23808 26056 23860
rect 26108 23848 26114 23860
rect 28445 23851 28503 23857
rect 28445 23848 28457 23851
rect 26108 23820 28457 23848
rect 26108 23808 26114 23820
rect 28445 23817 28457 23820
rect 28491 23817 28503 23851
rect 28445 23811 28503 23817
rect 28810 23808 28816 23860
rect 28868 23808 28874 23860
rect 14884 23752 15148 23780
rect 14884 23740 14890 23752
rect 8110 23672 8116 23724
rect 8168 23712 8174 23724
rect 13173 23715 13231 23721
rect 8168 23684 13124 23712
rect 8168 23672 8174 23684
rect 8846 23604 8852 23656
rect 8904 23644 8910 23656
rect 9582 23644 9588 23656
rect 8904 23616 9588 23644
rect 8904 23604 8910 23616
rect 9582 23604 9588 23616
rect 9640 23644 9646 23656
rect 12342 23644 12348 23656
rect 9640 23616 12348 23644
rect 9640 23604 9646 23616
rect 12342 23604 12348 23616
rect 12400 23604 12406 23656
rect 12713 23647 12771 23653
rect 12713 23613 12725 23647
rect 12759 23644 12771 23647
rect 12986 23644 12992 23656
rect 12759 23616 12992 23644
rect 12759 23613 12771 23616
rect 12713 23607 12771 23613
rect 12986 23604 12992 23616
rect 13044 23604 13050 23656
rect 13096 23576 13124 23684
rect 13173 23681 13185 23715
rect 13219 23681 13231 23715
rect 13173 23675 13231 23681
rect 13265 23715 13323 23721
rect 13265 23681 13277 23715
rect 13311 23712 13323 23715
rect 13906 23712 13912 23724
rect 13311 23684 13912 23712
rect 13311 23681 13323 23684
rect 13265 23675 13323 23681
rect 13188 23644 13216 23675
rect 13906 23672 13912 23684
rect 13964 23712 13970 23724
rect 14461 23715 14519 23721
rect 13964 23684 14412 23712
rect 13964 23672 13970 23684
rect 13538 23644 13544 23656
rect 13188 23616 13544 23644
rect 13538 23604 13544 23616
rect 13596 23644 13602 23656
rect 13814 23644 13820 23656
rect 13596 23616 13820 23644
rect 13596 23604 13602 23616
rect 13814 23604 13820 23616
rect 13872 23644 13878 23656
rect 14001 23647 14059 23653
rect 14001 23644 14013 23647
rect 13872 23616 14013 23644
rect 13872 23604 13878 23616
rect 14001 23613 14013 23616
rect 14047 23613 14059 23647
rect 14001 23607 14059 23613
rect 14090 23604 14096 23656
rect 14148 23604 14154 23656
rect 14384 23644 14412 23684
rect 14461 23681 14473 23715
rect 14507 23712 14519 23715
rect 14734 23712 14740 23724
rect 14507 23684 14740 23712
rect 14507 23681 14519 23684
rect 14461 23675 14519 23681
rect 14734 23672 14740 23684
rect 14792 23672 14798 23724
rect 15120 23721 15148 23752
rect 15565 23783 15623 23789
rect 15565 23749 15577 23783
rect 15611 23749 15623 23783
rect 15565 23743 15623 23749
rect 19610 23740 19616 23792
rect 19668 23740 19674 23792
rect 19702 23740 19708 23792
rect 19760 23780 19766 23792
rect 20257 23783 20315 23789
rect 19760 23752 20208 23780
rect 19760 23740 19766 23752
rect 15105 23715 15163 23721
rect 15105 23681 15117 23715
rect 15151 23681 15163 23715
rect 15105 23675 15163 23681
rect 15286 23672 15292 23724
rect 15344 23672 15350 23724
rect 15749 23715 15807 23721
rect 15749 23681 15761 23715
rect 15795 23681 15807 23715
rect 15749 23675 15807 23681
rect 19429 23715 19487 23721
rect 19429 23681 19441 23715
rect 19475 23712 19487 23715
rect 19720 23712 19748 23740
rect 19475 23684 19748 23712
rect 19475 23681 19487 23684
rect 19429 23675 19487 23681
rect 14826 23644 14832 23656
rect 14384 23616 14832 23644
rect 14826 23604 14832 23616
rect 14884 23644 14890 23656
rect 15013 23647 15071 23653
rect 15013 23644 15025 23647
rect 14884 23616 15025 23644
rect 14884 23604 14890 23616
rect 15013 23613 15025 23616
rect 15059 23613 15071 23647
rect 15764 23644 15792 23675
rect 19886 23672 19892 23724
rect 19944 23712 19950 23724
rect 20180 23721 20208 23752
rect 20257 23749 20269 23783
rect 20303 23780 20315 23783
rect 20438 23780 20444 23792
rect 20303 23752 20444 23780
rect 20303 23749 20315 23752
rect 20257 23743 20315 23749
rect 20438 23740 20444 23752
rect 20496 23780 20502 23792
rect 20625 23783 20683 23789
rect 20625 23780 20637 23783
rect 20496 23752 20637 23780
rect 20496 23740 20502 23752
rect 20625 23749 20637 23752
rect 20671 23749 20683 23783
rect 20732 23780 20760 23808
rect 24765 23783 24823 23789
rect 24765 23780 24777 23783
rect 20732 23752 24777 23780
rect 20625 23743 20683 23749
rect 20073 23715 20131 23721
rect 20073 23712 20085 23715
rect 19944 23684 20085 23712
rect 19944 23672 19950 23684
rect 20073 23681 20085 23684
rect 20119 23681 20131 23715
rect 20073 23675 20131 23681
rect 20165 23715 20223 23721
rect 20165 23681 20177 23715
rect 20211 23712 20223 23715
rect 20346 23712 20352 23724
rect 20211 23684 20352 23712
rect 20211 23681 20223 23684
rect 20165 23675 20223 23681
rect 20346 23672 20352 23684
rect 20404 23672 20410 23724
rect 21085 23715 21143 23721
rect 21085 23681 21097 23715
rect 21131 23681 21143 23715
rect 21085 23675 21143 23681
rect 15013 23607 15071 23613
rect 15212 23616 15792 23644
rect 14108 23576 14136 23604
rect 13096 23548 14136 23576
rect 9858 23468 9864 23520
rect 9916 23508 9922 23520
rect 10042 23508 10048 23520
rect 9916 23480 10048 23508
rect 9916 23468 9922 23480
rect 10042 23468 10048 23480
rect 10100 23468 10106 23520
rect 15010 23468 15016 23520
rect 15068 23508 15074 23520
rect 15212 23517 15240 23616
rect 19702 23604 19708 23656
rect 19760 23604 19766 23656
rect 20717 23647 20775 23653
rect 20717 23613 20729 23647
rect 20763 23644 20775 23647
rect 20990 23644 20996 23656
rect 20763 23616 20996 23644
rect 20763 23613 20775 23616
rect 20717 23607 20775 23613
rect 20990 23604 20996 23616
rect 21048 23604 21054 23656
rect 21100 23644 21128 23675
rect 21174 23672 21180 23724
rect 21232 23672 21238 23724
rect 23216 23721 23244 23752
rect 24765 23749 24777 23752
rect 24811 23749 24823 23783
rect 24765 23743 24823 23749
rect 27614 23740 27620 23792
rect 27672 23780 27678 23792
rect 28828 23780 28856 23808
rect 27672 23752 30604 23780
rect 27672 23740 27678 23752
rect 23201 23715 23259 23721
rect 23201 23681 23213 23715
rect 23247 23681 23259 23715
rect 23201 23675 23259 23681
rect 26418 23672 26424 23724
rect 26476 23672 26482 23724
rect 28074 23672 28080 23724
rect 28132 23712 28138 23724
rect 28353 23715 28411 23721
rect 28353 23712 28365 23715
rect 28132 23684 28365 23712
rect 28132 23672 28138 23684
rect 28353 23681 28365 23684
rect 28399 23681 28411 23715
rect 28353 23675 28411 23681
rect 28624 23715 28682 23721
rect 28624 23681 28636 23715
rect 28670 23681 28682 23715
rect 28624 23675 28682 23681
rect 21450 23644 21456 23656
rect 21100 23616 21456 23644
rect 21100 23588 21128 23616
rect 21450 23604 21456 23616
rect 21508 23604 21514 23656
rect 21634 23604 21640 23656
rect 21692 23604 21698 23656
rect 23477 23647 23535 23653
rect 23477 23613 23489 23647
rect 23523 23644 23535 23647
rect 23566 23644 23572 23656
rect 23523 23616 23572 23644
rect 23523 23613 23535 23616
rect 23477 23607 23535 23613
rect 23566 23604 23572 23616
rect 23624 23604 23630 23656
rect 27706 23604 27712 23656
rect 27764 23644 27770 23656
rect 27985 23647 28043 23653
rect 27985 23644 27997 23647
rect 27764 23616 27997 23644
rect 27764 23604 27770 23616
rect 27985 23613 27997 23616
rect 28031 23613 28043 23647
rect 27985 23607 28043 23613
rect 18230 23536 18236 23588
rect 18288 23576 18294 23588
rect 18874 23576 18880 23588
rect 18288 23548 18880 23576
rect 18288 23536 18294 23548
rect 18874 23536 18880 23548
rect 18932 23576 18938 23588
rect 19518 23576 19524 23588
rect 18932 23548 19524 23576
rect 18932 23536 18938 23548
rect 19518 23536 19524 23548
rect 19576 23576 19582 23588
rect 21082 23576 21088 23588
rect 19576 23548 21088 23576
rect 19576 23536 19582 23548
rect 21082 23536 21088 23548
rect 21140 23536 21146 23588
rect 24949 23579 25007 23585
rect 24949 23545 24961 23579
rect 24995 23576 25007 23579
rect 26694 23576 26700 23588
rect 24995 23548 26700 23576
rect 24995 23545 25007 23548
rect 24949 23539 25007 23545
rect 26694 23536 26700 23548
rect 26752 23536 26758 23588
rect 15197 23511 15255 23517
rect 15197 23508 15209 23511
rect 15068 23480 15209 23508
rect 15068 23468 15074 23480
rect 15197 23477 15209 23480
rect 15243 23477 15255 23511
rect 15197 23471 15255 23477
rect 15470 23468 15476 23520
rect 15528 23468 15534 23520
rect 26234 23468 26240 23520
rect 26292 23468 26298 23520
rect 27430 23468 27436 23520
rect 27488 23468 27494 23520
rect 27982 23468 27988 23520
rect 28040 23508 28046 23520
rect 28169 23511 28227 23517
rect 28169 23508 28181 23511
rect 28040 23480 28181 23508
rect 28040 23468 28046 23480
rect 28169 23477 28181 23480
rect 28215 23477 28227 23511
rect 28644 23508 28672 23675
rect 28718 23672 28724 23724
rect 28776 23672 28782 23724
rect 28810 23672 28816 23724
rect 28868 23672 28874 23724
rect 28996 23715 29054 23721
rect 28996 23681 29008 23715
rect 29042 23681 29054 23715
rect 28996 23675 29054 23681
rect 29089 23715 29147 23721
rect 29089 23681 29101 23715
rect 29135 23712 29147 23715
rect 29362 23712 29368 23724
rect 29135 23684 29368 23712
rect 29135 23681 29147 23684
rect 29089 23675 29147 23681
rect 28736 23576 28764 23672
rect 29012 23644 29040 23675
rect 29362 23672 29368 23684
rect 29420 23672 29426 23724
rect 30282 23672 30288 23724
rect 30340 23721 30346 23724
rect 30576 23721 30604 23752
rect 30340 23712 30352 23721
rect 30561 23715 30619 23721
rect 30340 23684 30385 23712
rect 30340 23675 30352 23684
rect 30561 23681 30573 23715
rect 30607 23681 30619 23715
rect 30561 23675 30619 23681
rect 30340 23672 30346 23675
rect 29546 23644 29552 23656
rect 29012 23616 29552 23644
rect 29546 23604 29552 23616
rect 29604 23604 29610 23656
rect 29181 23579 29239 23585
rect 29181 23576 29193 23579
rect 28736 23548 29193 23576
rect 29181 23545 29193 23548
rect 29227 23545 29239 23579
rect 29181 23539 29239 23545
rect 28718 23508 28724 23520
rect 28644 23480 28724 23508
rect 28169 23471 28227 23477
rect 28718 23468 28724 23480
rect 28776 23468 28782 23520
rect 1104 23418 31832 23440
rect 1104 23366 4182 23418
rect 4234 23366 4246 23418
rect 4298 23366 4310 23418
rect 4362 23366 4374 23418
rect 4426 23366 4438 23418
rect 4490 23366 4502 23418
rect 4554 23366 10182 23418
rect 10234 23366 10246 23418
rect 10298 23366 10310 23418
rect 10362 23366 10374 23418
rect 10426 23366 10438 23418
rect 10490 23366 10502 23418
rect 10554 23366 16182 23418
rect 16234 23366 16246 23418
rect 16298 23366 16310 23418
rect 16362 23366 16374 23418
rect 16426 23366 16438 23418
rect 16490 23366 16502 23418
rect 16554 23366 22182 23418
rect 22234 23366 22246 23418
rect 22298 23366 22310 23418
rect 22362 23366 22374 23418
rect 22426 23366 22438 23418
rect 22490 23366 22502 23418
rect 22554 23366 28182 23418
rect 28234 23366 28246 23418
rect 28298 23366 28310 23418
rect 28362 23366 28374 23418
rect 28426 23366 28438 23418
rect 28490 23366 28502 23418
rect 28554 23366 31832 23418
rect 1104 23344 31832 23366
rect 9398 23264 9404 23316
rect 9456 23304 9462 23316
rect 9456 23276 17632 23304
rect 9456 23264 9462 23276
rect 13906 23236 13912 23248
rect 6196 23208 13032 23236
rect 4157 23103 4215 23109
rect 4157 23069 4169 23103
rect 4203 23100 4215 23103
rect 4706 23100 4712 23112
rect 4203 23072 4712 23100
rect 4203 23069 4215 23072
rect 4157 23063 4215 23069
rect 4706 23060 4712 23072
rect 4764 23060 4770 23112
rect 5813 23103 5871 23109
rect 5813 23100 5825 23103
rect 4816 23072 5825 23100
rect 4816 22976 4844 23072
rect 5813 23069 5825 23072
rect 5859 23100 5871 23103
rect 5997 23103 6055 23109
rect 5997 23100 6009 23103
rect 5859 23072 6009 23100
rect 5859 23069 5871 23072
rect 5813 23063 5871 23069
rect 5997 23069 6009 23072
rect 6043 23069 6055 23103
rect 5997 23063 6055 23069
rect 5718 22992 5724 23044
rect 5776 23032 5782 23044
rect 6196 23041 6224 23208
rect 13004 23177 13032 23208
rect 13096 23208 13912 23236
rect 12989 23171 13047 23177
rect 12989 23137 13001 23171
rect 13035 23137 13047 23171
rect 12989 23131 13047 23137
rect 6365 23103 6423 23109
rect 6365 23069 6377 23103
rect 6411 23069 6423 23103
rect 6365 23063 6423 23069
rect 6181 23035 6239 23041
rect 6181 23032 6193 23035
rect 5776 23004 6193 23032
rect 5776 22992 5782 23004
rect 6181 23001 6193 23004
rect 6227 23001 6239 23035
rect 6181 22995 6239 23001
rect 6270 22992 6276 23044
rect 6328 22992 6334 23044
rect 6380 23032 6408 23063
rect 7926 23060 7932 23112
rect 7984 23100 7990 23112
rect 9493 23103 9551 23109
rect 9493 23100 9505 23103
rect 7984 23072 9505 23100
rect 7984 23060 7990 23072
rect 9493 23069 9505 23072
rect 9539 23069 9551 23103
rect 9493 23063 9551 23069
rect 12897 23103 12955 23109
rect 12897 23069 12909 23103
rect 12943 23100 12955 23103
rect 13096 23100 13124 23208
rect 13906 23196 13912 23208
rect 13964 23236 13970 23248
rect 14231 23239 14289 23245
rect 14231 23236 14243 23239
rect 13964 23208 14243 23236
rect 13964 23196 13970 23208
rect 14231 23205 14243 23208
rect 14277 23205 14289 23239
rect 14231 23199 14289 23205
rect 14369 23239 14427 23245
rect 14369 23205 14381 23239
rect 14415 23236 14427 23239
rect 14734 23236 14740 23248
rect 14415 23208 14740 23236
rect 14415 23205 14427 23208
rect 14369 23199 14427 23205
rect 14734 23196 14740 23208
rect 14792 23196 14798 23248
rect 15105 23239 15163 23245
rect 15105 23205 15117 23239
rect 15151 23236 15163 23239
rect 15930 23236 15936 23248
rect 15151 23208 15936 23236
rect 15151 23205 15163 23208
rect 15105 23199 15163 23205
rect 15930 23196 15936 23208
rect 15988 23196 15994 23248
rect 17604 23236 17632 23276
rect 18414 23264 18420 23316
rect 18472 23304 18478 23316
rect 19426 23304 19432 23316
rect 18472 23276 19432 23304
rect 18472 23264 18478 23276
rect 19426 23264 19432 23276
rect 19484 23264 19490 23316
rect 21542 23264 21548 23316
rect 21600 23304 21606 23316
rect 24118 23304 24124 23316
rect 21600 23276 24124 23304
rect 21600 23264 21606 23276
rect 24118 23264 24124 23276
rect 24176 23264 24182 23316
rect 27341 23307 27399 23313
rect 27341 23273 27353 23307
rect 27387 23304 27399 23307
rect 27706 23304 27712 23316
rect 27387 23276 27712 23304
rect 27387 23273 27399 23276
rect 27341 23267 27399 23273
rect 27706 23264 27712 23276
rect 27764 23264 27770 23316
rect 24854 23236 24860 23248
rect 17604 23208 24860 23236
rect 24854 23196 24860 23208
rect 24912 23196 24918 23248
rect 13814 23168 13820 23180
rect 13464 23140 13820 23168
rect 13464 23109 13492 23140
rect 13814 23128 13820 23140
rect 13872 23168 13878 23180
rect 14461 23171 14519 23177
rect 14461 23168 14473 23171
rect 13872 23140 14473 23168
rect 13872 23128 13878 23140
rect 14461 23137 14473 23140
rect 14507 23168 14519 23171
rect 14826 23168 14832 23180
rect 14507 23140 14832 23168
rect 14507 23137 14519 23140
rect 14461 23131 14519 23137
rect 14826 23128 14832 23140
rect 14884 23168 14890 23180
rect 19429 23171 19487 23177
rect 19429 23168 19441 23171
rect 14884 23140 19441 23168
rect 14884 23128 14890 23140
rect 12943 23072 13124 23100
rect 13357 23103 13415 23109
rect 12943 23069 12955 23072
rect 12897 23063 12955 23069
rect 13357 23069 13369 23103
rect 13403 23069 13415 23103
rect 13357 23063 13415 23069
rect 13449 23103 13507 23109
rect 13449 23069 13461 23103
rect 13495 23069 13507 23103
rect 13449 23063 13507 23069
rect 9858 23032 9864 23044
rect 6380 23004 9864 23032
rect 3973 22967 4031 22973
rect 3973 22933 3985 22967
rect 4019 22964 4031 22967
rect 4062 22964 4068 22976
rect 4019 22936 4068 22964
rect 4019 22933 4031 22936
rect 3973 22927 4031 22933
rect 4062 22924 4068 22936
rect 4120 22924 4126 22976
rect 4798 22924 4804 22976
rect 4856 22924 4862 22976
rect 5261 22967 5319 22973
rect 5261 22933 5273 22967
rect 5307 22964 5319 22967
rect 5442 22964 5448 22976
rect 5307 22936 5448 22964
rect 5307 22933 5319 22936
rect 5261 22927 5319 22933
rect 5442 22924 5448 22936
rect 5500 22924 5506 22976
rect 5902 22924 5908 22976
rect 5960 22964 5966 22976
rect 6380 22964 6408 23004
rect 9858 22992 9864 23004
rect 9916 22992 9922 23044
rect 12986 22992 12992 23044
rect 13044 23032 13050 23044
rect 13372 23032 13400 23063
rect 14366 23060 14372 23112
rect 14424 23100 14430 23112
rect 14921 23103 14979 23109
rect 14921 23100 14933 23103
rect 14424 23072 14933 23100
rect 14424 23060 14430 23072
rect 14921 23069 14933 23072
rect 14967 23069 14979 23103
rect 14921 23063 14979 23069
rect 15010 23060 15016 23112
rect 15068 23100 15074 23112
rect 15304 23109 15332 23140
rect 19429 23137 19441 23140
rect 19475 23168 19487 23171
rect 19794 23168 19800 23180
rect 19475 23140 19800 23168
rect 19475 23137 19487 23140
rect 19429 23131 19487 23137
rect 15105 23103 15163 23109
rect 15105 23100 15117 23103
rect 15068 23072 15117 23100
rect 15068 23060 15074 23072
rect 15105 23069 15117 23072
rect 15151 23069 15163 23103
rect 15105 23063 15163 23069
rect 15289 23103 15347 23109
rect 15289 23069 15301 23103
rect 15335 23069 15347 23103
rect 15289 23063 15347 23069
rect 15470 23060 15476 23112
rect 15528 23060 15534 23112
rect 15657 23103 15715 23109
rect 15657 23069 15669 23103
rect 15703 23069 15715 23103
rect 15657 23063 15715 23069
rect 13044 23004 13400 23032
rect 13541 23035 13599 23041
rect 13044 22992 13050 23004
rect 13541 23001 13553 23035
rect 13587 23032 13599 23035
rect 13630 23032 13636 23044
rect 13587 23004 13636 23032
rect 13587 23001 13599 23004
rect 13541 22995 13599 23001
rect 13630 22992 13636 23004
rect 13688 23032 13694 23044
rect 14090 23032 14096 23044
rect 13688 23004 14096 23032
rect 13688 22992 13694 23004
rect 14090 22992 14096 23004
rect 14148 22992 14154 23044
rect 15562 23032 15568 23044
rect 14292 23004 15568 23032
rect 5960 22936 6408 22964
rect 6549 22967 6607 22973
rect 5960 22924 5966 22936
rect 6549 22933 6561 22967
rect 6595 22964 6607 22967
rect 7742 22964 7748 22976
rect 6595 22936 7748 22964
rect 6595 22933 6607 22936
rect 6549 22927 6607 22933
rect 7742 22924 7748 22936
rect 7800 22924 7806 22976
rect 8938 22924 8944 22976
rect 8996 22924 9002 22976
rect 12802 22924 12808 22976
rect 12860 22964 12866 22976
rect 14292 22964 14320 23004
rect 15562 22992 15568 23004
rect 15620 22992 15626 23044
rect 15672 23032 15700 23063
rect 15746 23060 15752 23112
rect 15804 23100 15810 23112
rect 16301 23103 16359 23109
rect 16301 23100 16313 23103
rect 15804 23072 16313 23100
rect 15804 23060 15810 23072
rect 16301 23069 16313 23072
rect 16347 23069 16359 23103
rect 16301 23063 16359 23069
rect 18230 23060 18236 23112
rect 18288 23100 18294 23112
rect 18325 23103 18383 23109
rect 18325 23100 18337 23103
rect 18288 23072 18337 23100
rect 18288 23060 18294 23072
rect 18325 23069 18337 23072
rect 18371 23069 18383 23103
rect 18325 23063 18383 23069
rect 18598 23060 18604 23112
rect 18656 23060 18662 23112
rect 18785 23103 18843 23109
rect 18785 23069 18797 23103
rect 18831 23100 18843 23103
rect 18874 23100 18880 23112
rect 18831 23072 18880 23100
rect 18831 23069 18843 23072
rect 18785 23063 18843 23069
rect 18874 23060 18880 23072
rect 18932 23060 18938 23112
rect 15672 23004 15976 23032
rect 12860 22936 14320 22964
rect 14737 22967 14795 22973
rect 12860 22924 12866 22936
rect 14737 22933 14749 22967
rect 14783 22964 14795 22967
rect 15194 22964 15200 22976
rect 14783 22936 15200 22964
rect 14783 22933 14795 22936
rect 14737 22927 14795 22933
rect 15194 22924 15200 22936
rect 15252 22924 15258 22976
rect 15286 22924 15292 22976
rect 15344 22964 15350 22976
rect 15672 22964 15700 23004
rect 15344 22936 15700 22964
rect 15344 22924 15350 22936
rect 15838 22924 15844 22976
rect 15896 22924 15902 22976
rect 15948 22964 15976 23004
rect 16206 22992 16212 23044
rect 16264 23032 16270 23044
rect 16577 23035 16635 23041
rect 16577 23032 16589 23035
rect 16264 23004 16589 23032
rect 16264 22992 16270 23004
rect 16577 23001 16589 23004
rect 16623 23001 16635 23035
rect 16577 22995 16635 23001
rect 17586 22992 17592 23044
rect 17644 22992 17650 23044
rect 18414 22992 18420 23044
rect 18472 22992 18478 23044
rect 18432 22964 18460 22992
rect 15948 22936 18460 22964
rect 18506 22924 18512 22976
rect 18564 22924 18570 22976
rect 18969 22967 19027 22973
rect 18969 22933 18981 22967
rect 19015 22964 19027 22967
rect 19444 22964 19472 23131
rect 19794 23128 19800 23140
rect 19852 23128 19858 23180
rect 20346 23168 20352 23180
rect 19996 23140 20352 23168
rect 19610 23060 19616 23112
rect 19668 23100 19674 23112
rect 19996 23109 20024 23140
rect 20346 23128 20352 23140
rect 20404 23168 20410 23180
rect 21634 23168 21640 23180
rect 20404 23140 21640 23168
rect 20404 23128 20410 23140
rect 19889 23103 19947 23109
rect 19889 23100 19901 23103
rect 19668 23072 19901 23100
rect 19668 23060 19674 23072
rect 19889 23069 19901 23072
rect 19935 23069 19947 23103
rect 19889 23063 19947 23069
rect 19981 23103 20039 23109
rect 19981 23069 19993 23103
rect 20027 23069 20039 23103
rect 19981 23063 20039 23069
rect 20070 23060 20076 23112
rect 20128 23100 20134 23112
rect 20441 23103 20499 23109
rect 20441 23100 20453 23103
rect 20128 23072 20453 23100
rect 20128 23060 20134 23072
rect 20441 23069 20453 23072
rect 20487 23100 20499 23103
rect 20625 23103 20683 23109
rect 20625 23100 20637 23103
rect 20487 23072 20637 23100
rect 20487 23069 20499 23072
rect 20441 23063 20499 23069
rect 20625 23069 20637 23072
rect 20671 23069 20683 23103
rect 20625 23063 20683 23069
rect 21082 23060 21088 23112
rect 21140 23060 21146 23112
rect 21192 23109 21220 23140
rect 21634 23128 21640 23140
rect 21692 23168 21698 23180
rect 21692 23140 22416 23168
rect 21692 23128 21698 23140
rect 22388 23109 22416 23140
rect 25314 23128 25320 23180
rect 25372 23168 25378 23180
rect 25961 23171 26019 23177
rect 25961 23168 25973 23171
rect 25372 23140 25973 23168
rect 25372 23128 25378 23140
rect 25961 23137 25973 23140
rect 26007 23137 26019 23171
rect 25961 23131 26019 23137
rect 21177 23103 21235 23109
rect 21177 23069 21189 23103
rect 21223 23069 21235 23103
rect 21821 23103 21879 23109
rect 21821 23100 21833 23103
rect 21177 23063 21235 23069
rect 21284 23072 21680 23100
rect 20349 23035 20407 23041
rect 20349 23001 20361 23035
rect 20395 23001 20407 23035
rect 20349 22995 20407 23001
rect 19015 22936 19472 22964
rect 20364 22964 20392 22995
rect 20622 22964 20628 22976
rect 20364 22936 20628 22964
rect 19015 22933 19027 22936
rect 18969 22927 19027 22933
rect 20622 22924 20628 22936
rect 20680 22924 20686 22976
rect 21100 22964 21128 23060
rect 21284 23044 21312 23072
rect 21266 22992 21272 23044
rect 21324 22992 21330 23044
rect 21542 22992 21548 23044
rect 21600 22992 21606 23044
rect 21652 23041 21680 23072
rect 21744 23072 21833 23100
rect 21637 23035 21695 23041
rect 21637 23001 21649 23035
rect 21683 23001 21695 23035
rect 21637 22995 21695 23001
rect 21744 22976 21772 23072
rect 21821 23069 21833 23072
rect 21867 23069 21879 23103
rect 21821 23063 21879 23069
rect 22373 23103 22431 23109
rect 22373 23069 22385 23103
rect 22419 23100 22431 23103
rect 22554 23100 22560 23112
rect 22419 23072 22560 23100
rect 22419 23069 22431 23072
rect 22373 23063 22431 23069
rect 22554 23060 22560 23072
rect 22612 23060 22618 23112
rect 22833 23103 22891 23109
rect 22833 23100 22845 23103
rect 22664 23072 22845 23100
rect 22664 23044 22692 23072
rect 22833 23069 22845 23072
rect 22879 23069 22891 23103
rect 22833 23063 22891 23069
rect 23658 23060 23664 23112
rect 23716 23060 23722 23112
rect 24762 23060 24768 23112
rect 24820 23060 24826 23112
rect 25976 23100 26004 23131
rect 26050 23100 26056 23112
rect 25976 23072 26056 23100
rect 26050 23060 26056 23072
rect 26108 23100 26114 23112
rect 27525 23103 27583 23109
rect 27525 23100 27537 23103
rect 26108 23072 27537 23100
rect 26108 23060 26114 23072
rect 27525 23069 27537 23072
rect 27571 23100 27583 23103
rect 27614 23100 27620 23112
rect 27571 23072 27620 23100
rect 27571 23069 27583 23072
rect 27525 23063 27583 23069
rect 27614 23060 27620 23072
rect 27672 23060 27678 23112
rect 22278 22992 22284 23044
rect 22336 22992 22342 23044
rect 22646 22992 22652 23044
rect 22704 22992 22710 23044
rect 22738 22992 22744 23044
rect 22796 22992 22802 23044
rect 26234 23041 26240 23044
rect 26228 22995 26240 23041
rect 26292 23032 26298 23044
rect 27792 23035 27850 23041
rect 26292 23004 26328 23032
rect 26234 22992 26240 22995
rect 26292 22992 26298 23004
rect 27792 23001 27804 23035
rect 27838 23032 27850 23035
rect 27982 23032 27988 23044
rect 27838 23004 27988 23032
rect 27838 23001 27850 23004
rect 27792 22995 27850 23001
rect 27982 22992 27988 23004
rect 28040 22992 28046 23044
rect 21726 22964 21732 22976
rect 21100 22936 21732 22964
rect 21726 22924 21732 22936
rect 21784 22924 21790 22976
rect 23474 22924 23480 22976
rect 23532 22924 23538 22976
rect 25406 22924 25412 22976
rect 25464 22924 25470 22976
rect 28350 22924 28356 22976
rect 28408 22964 28414 22976
rect 28905 22967 28963 22973
rect 28905 22964 28917 22967
rect 28408 22936 28917 22964
rect 28408 22924 28414 22936
rect 28905 22933 28917 22936
rect 28951 22933 28963 22967
rect 28905 22927 28963 22933
rect 1104 22874 31832 22896
rect 1104 22822 4922 22874
rect 4974 22822 4986 22874
rect 5038 22822 5050 22874
rect 5102 22822 5114 22874
rect 5166 22822 5178 22874
rect 5230 22822 5242 22874
rect 5294 22822 10922 22874
rect 10974 22822 10986 22874
rect 11038 22822 11050 22874
rect 11102 22822 11114 22874
rect 11166 22822 11178 22874
rect 11230 22822 11242 22874
rect 11294 22822 16922 22874
rect 16974 22822 16986 22874
rect 17038 22822 17050 22874
rect 17102 22822 17114 22874
rect 17166 22822 17178 22874
rect 17230 22822 17242 22874
rect 17294 22822 22922 22874
rect 22974 22822 22986 22874
rect 23038 22822 23050 22874
rect 23102 22822 23114 22874
rect 23166 22822 23178 22874
rect 23230 22822 23242 22874
rect 23294 22822 28922 22874
rect 28974 22822 28986 22874
rect 29038 22822 29050 22874
rect 29102 22822 29114 22874
rect 29166 22822 29178 22874
rect 29230 22822 29242 22874
rect 29294 22822 31832 22874
rect 1104 22800 31832 22822
rect 3513 22763 3571 22769
rect 3513 22729 3525 22763
rect 3559 22729 3571 22763
rect 3513 22723 3571 22729
rect 3528 22692 3556 22723
rect 4798 22720 4804 22772
rect 4856 22760 4862 22772
rect 4985 22763 5043 22769
rect 4985 22760 4997 22763
rect 4856 22732 4997 22760
rect 4856 22720 4862 22732
rect 4985 22729 4997 22732
rect 5031 22729 5043 22763
rect 4985 22723 5043 22729
rect 5442 22720 5448 22772
rect 5500 22720 5506 22772
rect 7926 22720 7932 22772
rect 7984 22720 7990 22772
rect 8389 22763 8447 22769
rect 8389 22729 8401 22763
rect 8435 22760 8447 22763
rect 8938 22760 8944 22772
rect 8435 22732 8944 22760
rect 8435 22729 8447 22732
rect 8389 22723 8447 22729
rect 8938 22720 8944 22732
rect 8996 22720 9002 22772
rect 9858 22720 9864 22772
rect 9916 22720 9922 22772
rect 13814 22720 13820 22772
rect 13872 22720 13878 22772
rect 14366 22720 14372 22772
rect 14424 22760 14430 22772
rect 14553 22763 14611 22769
rect 14553 22760 14565 22763
rect 14424 22732 14565 22760
rect 14424 22720 14430 22732
rect 14553 22729 14565 22732
rect 14599 22729 14611 22763
rect 14553 22723 14611 22729
rect 15562 22720 15568 22772
rect 15620 22720 15626 22772
rect 15838 22720 15844 22772
rect 15896 22760 15902 22772
rect 16206 22760 16212 22772
rect 15896 22732 16212 22760
rect 15896 22720 15902 22732
rect 16206 22720 16212 22732
rect 16264 22720 16270 22772
rect 17954 22760 17960 22772
rect 16684 22732 17960 22760
rect 3850 22695 3908 22701
rect 3850 22692 3862 22695
rect 3528 22664 3862 22692
rect 3850 22661 3862 22664
rect 3896 22661 3908 22695
rect 3850 22655 3908 22661
rect 5350 22652 5356 22704
rect 5408 22692 5414 22704
rect 8662 22692 8668 22704
rect 5408 22664 8668 22692
rect 5408 22652 5414 22664
rect 6564 22633 6592 22664
rect 8662 22652 8668 22664
rect 8720 22652 8726 22704
rect 9876 22692 9904 22720
rect 12989 22695 13047 22701
rect 12989 22692 13001 22695
rect 9876 22664 13001 22692
rect 12989 22661 13001 22664
rect 13035 22661 13047 22695
rect 13832 22692 13860 22720
rect 12989 22655 13047 22661
rect 13372 22664 13860 22692
rect 3329 22627 3387 22633
rect 3329 22593 3341 22627
rect 3375 22593 3387 22627
rect 6549 22627 6607 22633
rect 3329 22587 3387 22593
rect 4632 22596 5672 22624
rect 3344 22420 3372 22587
rect 4632 22568 4660 22596
rect 3602 22516 3608 22568
rect 3660 22516 3666 22568
rect 4614 22516 4620 22568
rect 4672 22516 4678 22568
rect 5534 22516 5540 22568
rect 5592 22516 5598 22568
rect 5644 22565 5672 22596
rect 6549 22593 6561 22627
rect 6595 22593 6607 22627
rect 6549 22587 6607 22593
rect 6816 22627 6874 22633
rect 6816 22593 6828 22627
rect 6862 22624 6874 22627
rect 7282 22624 7288 22636
rect 6862 22596 7288 22624
rect 6862 22593 6874 22596
rect 6816 22587 6874 22593
rect 7282 22584 7288 22596
rect 7340 22584 7346 22636
rect 8481 22627 8539 22633
rect 8481 22593 8493 22627
rect 8527 22624 8539 22627
rect 9398 22624 9404 22636
rect 8527 22596 9404 22624
rect 8527 22593 8539 22596
rect 8481 22587 8539 22593
rect 9398 22584 9404 22596
rect 9456 22584 9462 22636
rect 13372 22633 13400 22664
rect 14090 22652 14096 22704
rect 14148 22692 14154 22704
rect 15580 22692 15608 22720
rect 14148 22664 14412 22692
rect 15580 22664 15792 22692
rect 14148 22652 14154 22664
rect 12897 22627 12955 22633
rect 12897 22593 12909 22627
rect 12943 22624 12955 22627
rect 13357 22627 13415 22633
rect 12943 22596 13032 22624
rect 12943 22593 12955 22596
rect 12897 22587 12955 22593
rect 13004 22568 13032 22596
rect 13357 22593 13369 22627
rect 13403 22593 13415 22627
rect 13357 22587 13415 22593
rect 13449 22627 13507 22633
rect 13449 22593 13461 22627
rect 13495 22593 13507 22627
rect 13449 22587 13507 22593
rect 13541 22627 13599 22633
rect 13541 22593 13553 22627
rect 13587 22624 13599 22627
rect 13906 22624 13912 22636
rect 13587 22596 13912 22624
rect 13587 22593 13599 22596
rect 13541 22587 13599 22593
rect 5629 22559 5687 22565
rect 5629 22525 5641 22559
rect 5675 22525 5687 22559
rect 5629 22519 5687 22525
rect 8570 22516 8576 22568
rect 8628 22556 8634 22568
rect 8665 22559 8723 22565
rect 8665 22556 8677 22559
rect 8628 22528 8677 22556
rect 8628 22516 8634 22528
rect 8665 22525 8677 22528
rect 8711 22556 8723 22559
rect 9582 22556 9588 22568
rect 8711 22528 9588 22556
rect 8711 22525 8723 22528
rect 8665 22519 8723 22525
rect 9582 22516 9588 22528
rect 9640 22516 9646 22568
rect 9858 22516 9864 22568
rect 9916 22556 9922 22568
rect 10042 22556 10048 22568
rect 9916 22528 10048 22556
rect 9916 22516 9922 22528
rect 10042 22516 10048 22528
rect 10100 22516 10106 22568
rect 12986 22516 12992 22568
rect 13044 22516 13050 22568
rect 13464 22556 13492 22587
rect 13906 22584 13912 22596
rect 13964 22624 13970 22636
rect 14384 22633 14412 22664
rect 14185 22627 14243 22633
rect 14185 22624 14197 22627
rect 13964 22596 14197 22624
rect 13964 22584 13970 22596
rect 14185 22593 14197 22596
rect 14231 22593 14243 22627
rect 14185 22587 14243 22593
rect 14369 22627 14427 22633
rect 14369 22593 14381 22627
rect 14415 22624 14427 22627
rect 14645 22627 14703 22633
rect 14645 22624 14657 22627
rect 14415 22596 14657 22624
rect 14415 22593 14427 22596
rect 14369 22587 14427 22593
rect 14645 22593 14657 22596
rect 14691 22624 14703 22627
rect 15562 22624 15568 22636
rect 14691 22596 15568 22624
rect 14691 22593 14703 22596
rect 14645 22587 14703 22593
rect 14090 22556 14096 22568
rect 13464 22528 14096 22556
rect 14090 22516 14096 22528
rect 14148 22516 14154 22568
rect 14200 22556 14228 22587
rect 15562 22584 15568 22596
rect 15620 22584 15626 22636
rect 15764 22633 15792 22664
rect 15749 22627 15807 22633
rect 15749 22593 15761 22627
rect 15795 22593 15807 22627
rect 15749 22587 15807 22593
rect 16022 22584 16028 22636
rect 16080 22624 16086 22636
rect 16684 22633 16712 22732
rect 17954 22720 17960 22732
rect 18012 22760 18018 22772
rect 18012 22732 20760 22760
rect 18012 22720 18018 22732
rect 18877 22695 18935 22701
rect 18877 22692 18889 22695
rect 18170 22664 18889 22692
rect 18877 22661 18889 22664
rect 18923 22661 18935 22695
rect 19334 22692 19340 22704
rect 18877 22655 18935 22661
rect 18984 22664 19340 22692
rect 18984 22633 19012 22664
rect 19334 22652 19340 22664
rect 19392 22692 19398 22704
rect 20732 22701 20760 22732
rect 20806 22720 20812 22772
rect 20864 22760 20870 22772
rect 20864 22732 23336 22760
rect 20864 22720 20870 22732
rect 19521 22695 19579 22701
rect 19521 22692 19533 22695
rect 19392 22664 19533 22692
rect 19392 22652 19398 22664
rect 19521 22661 19533 22664
rect 19567 22661 19579 22695
rect 20717 22695 20775 22701
rect 19521 22655 19579 22661
rect 19628 22664 20300 22692
rect 19628 22636 19656 22664
rect 16117 22627 16175 22633
rect 16117 22624 16129 22627
rect 16080 22596 16129 22624
rect 16080 22584 16086 22596
rect 16117 22593 16129 22596
rect 16163 22593 16175 22627
rect 16117 22587 16175 22593
rect 16669 22627 16727 22633
rect 16669 22593 16681 22627
rect 16715 22593 16727 22627
rect 18969 22627 19027 22633
rect 18969 22624 18981 22627
rect 16669 22587 16727 22593
rect 18616 22596 18981 22624
rect 15841 22559 15899 22565
rect 15841 22556 15853 22559
rect 14200 22528 15853 22556
rect 15841 22525 15853 22528
rect 15887 22525 15899 22559
rect 15841 22519 15899 22525
rect 5077 22491 5135 22497
rect 5077 22488 5089 22491
rect 4540 22460 5089 22488
rect 4540 22420 4568 22460
rect 5077 22457 5089 22460
rect 5123 22457 5135 22491
rect 15856 22488 15884 22519
rect 15930 22516 15936 22568
rect 15988 22516 15994 22568
rect 16301 22559 16359 22565
rect 16301 22525 16313 22559
rect 16347 22556 16359 22559
rect 16945 22559 17003 22565
rect 16945 22556 16957 22559
rect 16347 22528 16957 22556
rect 16347 22525 16359 22528
rect 16301 22519 16359 22525
rect 16945 22525 16957 22528
rect 16991 22525 17003 22559
rect 16945 22519 17003 22525
rect 18616 22500 18644 22596
rect 18969 22593 18981 22596
rect 19015 22593 19027 22627
rect 18969 22587 19027 22593
rect 19058 22584 19064 22636
rect 19116 22624 19122 22636
rect 19245 22627 19303 22633
rect 19245 22624 19257 22627
rect 19116 22596 19257 22624
rect 19116 22584 19122 22596
rect 19245 22593 19257 22596
rect 19291 22593 19303 22627
rect 19245 22587 19303 22593
rect 19610 22584 19616 22636
rect 19668 22584 19674 22636
rect 19797 22627 19855 22633
rect 19797 22593 19809 22627
rect 19843 22624 19855 22627
rect 19978 22624 19984 22636
rect 19843 22596 19984 22624
rect 19843 22593 19855 22596
rect 19797 22587 19855 22593
rect 18693 22559 18751 22565
rect 18693 22525 18705 22559
rect 18739 22556 18751 22559
rect 19812 22556 19840 22587
rect 19978 22584 19984 22596
rect 20036 22584 20042 22636
rect 20070 22584 20076 22636
rect 20128 22584 20134 22636
rect 20272 22633 20300 22664
rect 20717 22661 20729 22695
rect 20763 22692 20775 22695
rect 22830 22692 22836 22704
rect 20763 22664 22836 22692
rect 20763 22661 20775 22664
rect 20717 22655 20775 22661
rect 22830 22652 22836 22664
rect 22888 22692 22894 22704
rect 22888 22664 23152 22692
rect 22888 22652 22894 22664
rect 20257 22627 20315 22633
rect 20257 22593 20269 22627
rect 20303 22593 20315 22627
rect 20257 22587 20315 22593
rect 18739 22528 19840 22556
rect 18739 22525 18751 22528
rect 18693 22519 18751 22525
rect 5077 22451 5135 22457
rect 12406 22460 15240 22488
rect 15856 22460 15976 22488
rect 3344 22392 4568 22420
rect 8018 22380 8024 22432
rect 8076 22380 8082 22432
rect 11054 22380 11060 22432
rect 11112 22420 11118 22432
rect 12158 22420 12164 22432
rect 11112 22392 12164 22420
rect 11112 22380 11118 22392
rect 12158 22380 12164 22392
rect 12216 22420 12222 22432
rect 12406 22420 12434 22460
rect 15212 22432 15240 22460
rect 12216 22392 12434 22420
rect 14277 22423 14335 22429
rect 12216 22380 12222 22392
rect 14277 22389 14289 22423
rect 14323 22420 14335 22423
rect 14642 22420 14648 22432
rect 14323 22392 14648 22420
rect 14323 22389 14335 22392
rect 14277 22383 14335 22389
rect 14642 22380 14648 22392
rect 14700 22380 14706 22432
rect 15194 22380 15200 22432
rect 15252 22380 15258 22432
rect 15749 22423 15807 22429
rect 15749 22389 15761 22423
rect 15795 22420 15807 22423
rect 15838 22420 15844 22432
rect 15795 22392 15844 22420
rect 15795 22389 15807 22392
rect 15749 22383 15807 22389
rect 15838 22380 15844 22392
rect 15896 22380 15902 22432
rect 15948 22420 15976 22460
rect 18598 22448 18604 22500
rect 18656 22448 18662 22500
rect 19981 22491 20039 22497
rect 19981 22457 19993 22491
rect 20027 22488 20039 22491
rect 20088 22488 20116 22584
rect 20027 22460 20116 22488
rect 20272 22488 20300 22587
rect 20898 22584 20904 22636
rect 20956 22624 20962 22636
rect 21545 22627 21603 22633
rect 21545 22624 21557 22627
rect 20956 22596 21557 22624
rect 20956 22584 20962 22596
rect 21545 22593 21557 22596
rect 21591 22593 21603 22627
rect 21545 22587 21603 22593
rect 21726 22584 21732 22636
rect 21784 22624 21790 22636
rect 22465 22627 22523 22633
rect 22465 22624 22477 22627
rect 21784 22596 22477 22624
rect 21784 22584 21790 22596
rect 22465 22593 22477 22596
rect 22511 22593 22523 22627
rect 22465 22587 22523 22593
rect 22554 22584 22560 22636
rect 22612 22584 22618 22636
rect 22646 22584 22652 22636
rect 22704 22584 22710 22636
rect 23124 22633 23152 22664
rect 23109 22627 23167 22633
rect 23109 22593 23121 22627
rect 23155 22593 23167 22627
rect 23308 22624 23336 22732
rect 23474 22720 23480 22772
rect 23532 22720 23538 22772
rect 23658 22720 23664 22772
rect 23716 22760 23722 22772
rect 24581 22763 24639 22769
rect 24581 22760 24593 22763
rect 23716 22732 24593 22760
rect 23716 22720 23722 22732
rect 24581 22729 24593 22732
rect 24627 22729 24639 22763
rect 24581 22723 24639 22729
rect 24949 22763 25007 22769
rect 24949 22729 24961 22763
rect 24995 22760 25007 22763
rect 25406 22760 25412 22772
rect 24995 22732 25412 22760
rect 24995 22729 25007 22732
rect 24949 22723 25007 22729
rect 25406 22720 25412 22732
rect 25464 22720 25470 22772
rect 27706 22760 27712 22772
rect 26344 22732 27712 22760
rect 23376 22695 23434 22701
rect 23376 22661 23388 22695
rect 23422 22692 23434 22695
rect 23492 22692 23520 22720
rect 23422 22664 23520 22692
rect 23422 22661 23434 22664
rect 23376 22655 23434 22661
rect 23842 22652 23848 22704
rect 23900 22692 23906 22704
rect 25041 22695 25099 22701
rect 25041 22692 25053 22695
rect 23900 22664 25053 22692
rect 23900 22652 23906 22664
rect 25041 22661 25053 22664
rect 25087 22661 25099 22695
rect 25041 22655 25099 22661
rect 26257 22627 26315 22633
rect 23308 22596 25360 22624
rect 23109 22587 23167 22593
rect 21450 22516 21456 22568
rect 21508 22556 21514 22568
rect 22278 22556 22284 22568
rect 21508 22528 22284 22556
rect 21508 22516 21514 22528
rect 22278 22516 22284 22528
rect 22336 22556 22342 22568
rect 22373 22559 22431 22565
rect 22373 22556 22385 22559
rect 22336 22528 22385 22556
rect 22336 22516 22342 22528
rect 22373 22525 22385 22528
rect 22419 22525 22431 22559
rect 22373 22519 22431 22525
rect 22664 22488 22692 22584
rect 25222 22516 25228 22568
rect 25280 22516 25286 22568
rect 25332 22556 25360 22596
rect 26257 22593 26269 22627
rect 26303 22624 26315 22627
rect 26344 22624 26372 22732
rect 27706 22720 27712 22732
rect 27764 22720 27770 22772
rect 28074 22720 28080 22772
rect 28132 22760 28138 22772
rect 28445 22763 28503 22769
rect 28445 22760 28457 22763
rect 28132 22732 28457 22760
rect 28132 22720 28138 22732
rect 28445 22729 28457 22732
rect 28491 22729 28503 22763
rect 28445 22723 28503 22729
rect 28626 22720 28632 22772
rect 28684 22760 28690 22772
rect 28905 22763 28963 22769
rect 28905 22760 28917 22763
rect 28684 22732 28917 22760
rect 28684 22720 28690 22732
rect 28905 22729 28917 22732
rect 28951 22729 28963 22763
rect 28905 22723 28963 22729
rect 26421 22695 26479 22701
rect 26421 22661 26433 22695
rect 26467 22661 26479 22695
rect 26421 22655 26479 22661
rect 26513 22695 26571 22701
rect 26513 22661 26525 22695
rect 26559 22692 26571 22695
rect 28350 22692 28356 22704
rect 26559 22664 28356 22692
rect 26559 22661 26571 22664
rect 26513 22655 26571 22661
rect 26303 22596 26372 22624
rect 26303 22593 26315 22596
rect 26257 22587 26315 22593
rect 26436 22556 26464 22655
rect 28350 22652 28356 22664
rect 28408 22692 28414 22704
rect 28408 22664 29868 22692
rect 28408 22652 28414 22664
rect 26605 22627 26663 22633
rect 26605 22593 26617 22627
rect 26651 22624 26663 22627
rect 27154 22624 27160 22636
rect 26651 22596 27160 22624
rect 26651 22593 26663 22596
rect 26605 22587 26663 22593
rect 27154 22584 27160 22596
rect 27212 22584 27218 22636
rect 27338 22584 27344 22636
rect 27396 22584 27402 22636
rect 29840 22633 29868 22664
rect 27801 22627 27859 22633
rect 27801 22593 27813 22627
rect 27847 22624 27859 22627
rect 28813 22627 28871 22633
rect 27847 22596 28764 22624
rect 27847 22593 27859 22596
rect 27801 22587 27859 22593
rect 26878 22556 26884 22568
rect 25332 22528 26884 22556
rect 26878 22516 26884 22528
rect 26936 22556 26942 22568
rect 27356 22556 27384 22584
rect 28736 22568 28764 22596
rect 28813 22593 28825 22627
rect 28859 22624 28871 22627
rect 29273 22627 29331 22633
rect 29273 22624 29285 22627
rect 28859 22596 29285 22624
rect 28859 22593 28871 22596
rect 28813 22587 28871 22593
rect 29273 22593 29285 22596
rect 29319 22593 29331 22627
rect 29273 22587 29331 22593
rect 29825 22627 29883 22633
rect 29825 22593 29837 22627
rect 29871 22593 29883 22627
rect 29825 22587 29883 22593
rect 26936 22528 27384 22556
rect 27525 22559 27583 22565
rect 26936 22516 26942 22528
rect 27525 22525 27537 22559
rect 27571 22525 27583 22559
rect 27525 22519 27583 22525
rect 20272 22460 22692 22488
rect 22833 22491 22891 22497
rect 20027 22457 20039 22460
rect 19981 22451 20039 22457
rect 22833 22457 22845 22491
rect 22879 22457 22891 22491
rect 27540 22488 27568 22519
rect 28718 22516 28724 22568
rect 28776 22516 28782 22568
rect 28997 22559 29055 22565
rect 28997 22525 29009 22559
rect 29043 22525 29055 22559
rect 28997 22519 29055 22525
rect 22833 22451 22891 22457
rect 24412 22460 27568 22488
rect 19996 22420 20024 22451
rect 15948 22392 20024 22420
rect 20441 22423 20499 22429
rect 20441 22389 20453 22423
rect 20487 22420 20499 22423
rect 21266 22420 21272 22432
rect 20487 22392 21272 22420
rect 20487 22389 20499 22392
rect 20441 22383 20499 22389
rect 21266 22380 21272 22392
rect 21324 22380 21330 22432
rect 22848 22420 22876 22451
rect 24412 22420 24440 22460
rect 27982 22448 27988 22500
rect 28040 22488 28046 22500
rect 29012 22488 29040 22519
rect 28040 22460 29040 22488
rect 28040 22448 28046 22460
rect 22848 22392 24440 22420
rect 24489 22423 24547 22429
rect 24489 22389 24501 22423
rect 24535 22420 24547 22423
rect 24762 22420 24768 22432
rect 24535 22392 24768 22420
rect 24535 22389 24547 22392
rect 24489 22383 24547 22389
rect 24762 22380 24768 22392
rect 24820 22380 24826 22432
rect 26786 22380 26792 22432
rect 26844 22380 26850 22432
rect 1104 22330 31832 22352
rect 1104 22278 4182 22330
rect 4234 22278 4246 22330
rect 4298 22278 4310 22330
rect 4362 22278 4374 22330
rect 4426 22278 4438 22330
rect 4490 22278 4502 22330
rect 4554 22278 10182 22330
rect 10234 22278 10246 22330
rect 10298 22278 10310 22330
rect 10362 22278 10374 22330
rect 10426 22278 10438 22330
rect 10490 22278 10502 22330
rect 10554 22278 16182 22330
rect 16234 22278 16246 22330
rect 16298 22278 16310 22330
rect 16362 22278 16374 22330
rect 16426 22278 16438 22330
rect 16490 22278 16502 22330
rect 16554 22278 22182 22330
rect 22234 22278 22246 22330
rect 22298 22278 22310 22330
rect 22362 22278 22374 22330
rect 22426 22278 22438 22330
rect 22490 22278 22502 22330
rect 22554 22278 28182 22330
rect 28234 22278 28246 22330
rect 28298 22278 28310 22330
rect 28362 22278 28374 22330
rect 28426 22278 28438 22330
rect 28490 22278 28502 22330
rect 28554 22278 31832 22330
rect 1104 22256 31832 22278
rect 4706 22176 4712 22228
rect 4764 22216 4770 22228
rect 5261 22219 5319 22225
rect 5261 22216 5273 22219
rect 4764 22188 5273 22216
rect 4764 22176 4770 22188
rect 5261 22185 5273 22188
rect 5307 22185 5319 22219
rect 5261 22179 5319 22185
rect 7282 22176 7288 22228
rect 7340 22176 7346 22228
rect 8018 22176 8024 22228
rect 8076 22176 8082 22228
rect 10134 22176 10140 22228
rect 10192 22216 10198 22228
rect 10321 22219 10379 22225
rect 10321 22216 10333 22219
rect 10192 22188 10333 22216
rect 10192 22176 10198 22188
rect 10321 22185 10333 22188
rect 10367 22185 10379 22219
rect 10321 22179 10379 22185
rect 15856 22188 18276 22216
rect 5810 22108 5816 22160
rect 5868 22148 5874 22160
rect 5994 22148 6000 22160
rect 5868 22120 6000 22148
rect 5868 22108 5874 22120
rect 5920 22089 5948 22120
rect 5994 22108 6000 22120
rect 6052 22108 6058 22160
rect 5905 22083 5963 22089
rect 5905 22049 5917 22083
rect 5951 22080 5963 22083
rect 8036 22080 8064 22176
rect 9953 22151 10011 22157
rect 9953 22148 9965 22151
rect 9784 22120 9965 22148
rect 5951 22052 5985 22080
rect 7484 22052 8064 22080
rect 5951 22049 5963 22052
rect 5905 22043 5963 22049
rect 3602 21972 3608 22024
rect 3660 22012 3666 22024
rect 3789 22015 3847 22021
rect 3789 22012 3801 22015
rect 3660 21984 3801 22012
rect 3660 21972 3666 21984
rect 3789 21981 3801 21984
rect 3835 22012 3847 22015
rect 5350 22012 5356 22024
rect 3835 21984 5356 22012
rect 3835 21981 3847 21984
rect 3789 21975 3847 21981
rect 5350 21972 5356 21984
rect 5408 21972 5414 22024
rect 7484 22021 7512 22052
rect 9582 22040 9588 22092
rect 9640 22080 9646 22092
rect 9784 22080 9812 22120
rect 9953 22117 9965 22120
rect 9999 22117 10011 22151
rect 9953 22111 10011 22117
rect 10226 22108 10232 22160
rect 10284 22148 10290 22160
rect 10778 22148 10784 22160
rect 10284 22120 10784 22148
rect 10284 22108 10290 22120
rect 10778 22108 10784 22120
rect 10836 22148 10842 22160
rect 10836 22120 12664 22148
rect 10836 22108 10842 22120
rect 12636 22089 12664 22120
rect 15562 22108 15568 22160
rect 15620 22148 15626 22160
rect 15856 22148 15884 22188
rect 15620 22120 15884 22148
rect 18248 22148 18276 22188
rect 19978 22176 19984 22228
rect 20036 22216 20042 22228
rect 21450 22216 21456 22228
rect 20036 22188 21456 22216
rect 20036 22176 20042 22188
rect 21450 22176 21456 22188
rect 21508 22176 21514 22228
rect 21545 22219 21603 22225
rect 21545 22185 21557 22219
rect 21591 22216 21603 22219
rect 21634 22216 21640 22228
rect 21591 22188 21640 22216
rect 21591 22185 21603 22188
rect 21545 22179 21603 22185
rect 21634 22176 21640 22188
rect 21692 22176 21698 22228
rect 21266 22148 21272 22160
rect 18248 22120 21272 22148
rect 15620 22108 15626 22120
rect 21266 22108 21272 22120
rect 21324 22108 21330 22160
rect 24026 22108 24032 22160
rect 24084 22148 24090 22160
rect 24084 22120 24992 22148
rect 24084 22108 24090 22120
rect 10689 22083 10747 22089
rect 10689 22080 10701 22083
rect 9640 22052 9812 22080
rect 9876 22052 10701 22080
rect 9640 22040 9646 22052
rect 7193 22015 7251 22021
rect 7193 21981 7205 22015
rect 7239 21981 7251 22015
rect 7193 21975 7251 21981
rect 7469 22015 7527 22021
rect 7469 21981 7481 22015
rect 7515 21981 7527 22015
rect 7469 21975 7527 21981
rect 4062 21953 4068 21956
rect 4056 21907 4068 21953
rect 4062 21904 4068 21907
rect 4120 21904 4126 21956
rect 5184 21916 6316 21944
rect 5184 21885 5212 21916
rect 6288 21888 6316 21916
rect 7208 21888 7236 21975
rect 7742 21972 7748 22024
rect 7800 21972 7806 22024
rect 7926 21972 7932 22024
rect 7984 21972 7990 22024
rect 8018 21972 8024 22024
rect 8076 21972 8082 22024
rect 8205 22015 8263 22021
rect 8205 21981 8217 22015
rect 8251 22012 8263 22015
rect 8938 22012 8944 22024
rect 8251 21984 8944 22012
rect 8251 21981 8263 21984
rect 8205 21975 8263 21981
rect 8938 21972 8944 21984
rect 8996 21972 9002 22024
rect 9876 22021 9904 22052
rect 10689 22049 10701 22052
rect 10735 22049 10747 22083
rect 10689 22043 10747 22049
rect 12621 22083 12679 22089
rect 12621 22049 12633 22083
rect 12667 22080 12679 22083
rect 15746 22080 15752 22092
rect 12667 22052 15752 22080
rect 12667 22049 12679 22052
rect 12621 22043 12679 22049
rect 15746 22040 15752 22052
rect 15804 22040 15810 22092
rect 15838 22040 15844 22092
rect 15896 22080 15902 22092
rect 16945 22083 17003 22089
rect 15896 22052 16344 22080
rect 15896 22040 15902 22052
rect 9861 22015 9919 22021
rect 9861 21981 9873 22015
rect 9907 21981 9919 22015
rect 10045 22015 10103 22021
rect 10045 22012 10057 22015
rect 9861 21975 9919 21981
rect 9968 21984 10057 22012
rect 7561 21947 7619 21953
rect 7561 21913 7573 21947
rect 7607 21944 7619 21947
rect 7607 21916 8800 21944
rect 7607 21913 7619 21916
rect 7561 21907 7619 21913
rect 5169 21879 5227 21885
rect 5169 21845 5181 21879
rect 5215 21845 5227 21879
rect 5169 21839 5227 21845
rect 5626 21836 5632 21888
rect 5684 21836 5690 21888
rect 5721 21879 5779 21885
rect 5721 21845 5733 21879
rect 5767 21876 5779 21879
rect 6086 21876 6092 21888
rect 5767 21848 6092 21876
rect 5767 21845 5779 21848
rect 5721 21839 5779 21845
rect 6086 21836 6092 21848
rect 6144 21836 6150 21888
rect 6270 21836 6276 21888
rect 6328 21836 6334 21888
rect 6546 21836 6552 21888
rect 6604 21836 6610 21888
rect 7190 21836 7196 21888
rect 7248 21836 7254 21888
rect 8389 21879 8447 21885
rect 8389 21845 8401 21879
rect 8435 21876 8447 21879
rect 8478 21876 8484 21888
rect 8435 21848 8484 21876
rect 8435 21845 8447 21848
rect 8389 21839 8447 21845
rect 8478 21836 8484 21848
rect 8536 21836 8542 21888
rect 8772 21876 8800 21916
rect 9214 21904 9220 21956
rect 9272 21944 9278 21956
rect 9398 21944 9404 21956
rect 9272 21916 9404 21944
rect 9272 21904 9278 21916
rect 9398 21904 9404 21916
rect 9456 21904 9462 21956
rect 9968 21876 9996 21984
rect 10045 21981 10057 21984
rect 10091 21981 10103 22015
rect 10045 21975 10103 21981
rect 10137 22015 10195 22021
rect 10137 21981 10149 22015
rect 10183 22012 10195 22015
rect 10183 21984 10548 22012
rect 10183 21981 10195 21984
rect 10137 21975 10195 21981
rect 8772 21848 9996 21876
rect 10410 21836 10416 21888
rect 10468 21836 10474 21888
rect 10520 21876 10548 21984
rect 10594 21972 10600 22024
rect 10652 21972 10658 22024
rect 11054 21972 11060 22024
rect 11112 21972 11118 22024
rect 16114 21972 16120 22024
rect 16172 21972 16178 22024
rect 16316 22021 16344 22052
rect 16945 22049 16957 22083
rect 16991 22080 17003 22083
rect 16991 22052 20024 22080
rect 16991 22049 17003 22052
rect 16945 22043 17003 22049
rect 16301 22015 16359 22021
rect 16301 21981 16313 22015
rect 16347 21981 16359 22015
rect 18506 22012 18512 22024
rect 18354 21984 18512 22012
rect 16301 21975 16359 21981
rect 18506 21972 18512 21984
rect 18564 21972 18570 22024
rect 18969 22015 19027 22021
rect 18969 21981 18981 22015
rect 19015 22012 19027 22015
rect 19610 22012 19616 22024
rect 19015 21984 19616 22012
rect 19015 21981 19027 21984
rect 18969 21975 19027 21981
rect 19610 21972 19616 21984
rect 19668 21972 19674 22024
rect 19996 21956 20024 22052
rect 21284 22021 21312 22108
rect 21637 22083 21695 22089
rect 21637 22049 21649 22083
rect 21683 22080 21695 22083
rect 21726 22080 21732 22092
rect 21683 22052 21732 22080
rect 21683 22049 21695 22052
rect 21637 22043 21695 22049
rect 21726 22040 21732 22052
rect 21784 22040 21790 22092
rect 22830 22040 22836 22092
rect 22888 22040 22894 22092
rect 24854 22040 24860 22092
rect 24912 22040 24918 22092
rect 24964 22089 24992 22120
rect 24949 22083 25007 22089
rect 24949 22049 24961 22083
rect 24995 22080 25007 22083
rect 24995 22052 25029 22080
rect 24995 22049 25007 22052
rect 24949 22043 25007 22049
rect 26418 22040 26424 22092
rect 26476 22040 26482 22092
rect 27522 22040 27528 22092
rect 27580 22040 27586 22092
rect 21269 22015 21327 22021
rect 21269 21981 21281 22015
rect 21315 21981 21327 22015
rect 26436 22012 26464 22040
rect 27341 22015 27399 22021
rect 21269 21975 21327 21981
rect 22066 21984 24992 22012
rect 26436 21984 26740 22012
rect 10778 21904 10784 21956
rect 10836 21944 10842 21956
rect 10873 21947 10931 21953
rect 10873 21944 10885 21947
rect 10836 21916 10885 21944
rect 10836 21904 10842 21916
rect 10873 21913 10885 21916
rect 10919 21913 10931 21947
rect 10873 21907 10931 21913
rect 11330 21904 11336 21956
rect 11388 21944 11394 21956
rect 11793 21947 11851 21953
rect 11793 21944 11805 21947
rect 11388 21916 11805 21944
rect 11388 21904 11394 21916
rect 11793 21913 11805 21916
rect 11839 21913 11851 21947
rect 11793 21907 11851 21913
rect 16209 21947 16267 21953
rect 16209 21913 16221 21947
rect 16255 21944 16267 21947
rect 17221 21947 17279 21953
rect 17221 21944 17233 21947
rect 16255 21916 17233 21944
rect 16255 21913 16267 21916
rect 16209 21907 16267 21913
rect 17221 21913 17233 21916
rect 17267 21913 17279 21947
rect 17221 21907 17279 21913
rect 19978 21904 19984 21956
rect 20036 21904 20042 21956
rect 20714 21904 20720 21956
rect 20772 21904 20778 21956
rect 17310 21876 17316 21888
rect 10520 21848 17316 21876
rect 17310 21836 17316 21848
rect 17368 21836 17374 21888
rect 21361 21879 21419 21885
rect 21361 21845 21373 21879
rect 21407 21876 21419 21879
rect 22066 21876 22094 21984
rect 23100 21947 23158 21953
rect 23100 21913 23112 21947
rect 23146 21944 23158 21947
rect 23474 21944 23480 21956
rect 23146 21916 23480 21944
rect 23146 21913 23158 21916
rect 23100 21907 23158 21913
rect 23474 21904 23480 21916
rect 23532 21904 23538 21956
rect 23676 21916 24440 21944
rect 23676 21888 23704 21916
rect 21407 21848 22094 21876
rect 21407 21845 21419 21848
rect 21361 21839 21419 21845
rect 23658 21836 23664 21888
rect 23716 21836 23722 21888
rect 24210 21836 24216 21888
rect 24268 21836 24274 21888
rect 24412 21885 24440 21916
rect 24397 21879 24455 21885
rect 24397 21845 24409 21879
rect 24443 21845 24455 21879
rect 24397 21839 24455 21845
rect 24762 21836 24768 21888
rect 24820 21836 24826 21888
rect 24964 21876 24992 21984
rect 25314 21904 25320 21956
rect 25372 21944 25378 21956
rect 25685 21947 25743 21953
rect 25685 21944 25697 21947
rect 25372 21916 25697 21944
rect 25372 21904 25378 21916
rect 25685 21913 25697 21916
rect 25731 21913 25743 21947
rect 25685 21907 25743 21913
rect 26142 21904 26148 21956
rect 26200 21944 26206 21956
rect 26421 21947 26479 21953
rect 26421 21944 26433 21947
rect 26200 21916 26433 21944
rect 26200 21904 26206 21916
rect 26421 21913 26433 21916
rect 26467 21913 26479 21947
rect 26421 21907 26479 21913
rect 26234 21876 26240 21888
rect 24964 21848 26240 21876
rect 26234 21836 26240 21848
rect 26292 21836 26298 21888
rect 26712 21876 26740 21984
rect 27341 21981 27353 22015
rect 27387 22012 27399 22015
rect 27430 22012 27436 22024
rect 27387 21984 27436 22012
rect 27387 21981 27399 21984
rect 27341 21975 27399 21981
rect 27430 21972 27436 21984
rect 27488 21972 27494 22024
rect 29638 21972 29644 22024
rect 29696 22012 29702 22024
rect 30101 22015 30159 22021
rect 30101 22012 30113 22015
rect 29696 21984 30113 22012
rect 29696 21972 29702 21984
rect 30101 21981 30113 21984
rect 30147 21981 30159 22015
rect 30101 21975 30159 21981
rect 26973 21879 27031 21885
rect 26973 21876 26985 21879
rect 26712 21848 26985 21876
rect 26973 21845 26985 21848
rect 27019 21845 27031 21879
rect 26973 21839 27031 21845
rect 27430 21836 27436 21888
rect 27488 21836 27494 21888
rect 29546 21836 29552 21888
rect 29604 21836 29610 21888
rect 1104 21786 31832 21808
rect 1104 21734 4922 21786
rect 4974 21734 4986 21786
rect 5038 21734 5050 21786
rect 5102 21734 5114 21786
rect 5166 21734 5178 21786
rect 5230 21734 5242 21786
rect 5294 21734 10922 21786
rect 10974 21734 10986 21786
rect 11038 21734 11050 21786
rect 11102 21734 11114 21786
rect 11166 21734 11178 21786
rect 11230 21734 11242 21786
rect 11294 21734 16922 21786
rect 16974 21734 16986 21786
rect 17038 21734 17050 21786
rect 17102 21734 17114 21786
rect 17166 21734 17178 21786
rect 17230 21734 17242 21786
rect 17294 21734 22922 21786
rect 22974 21734 22986 21786
rect 23038 21734 23050 21786
rect 23102 21734 23114 21786
rect 23166 21734 23178 21786
rect 23230 21734 23242 21786
rect 23294 21734 28922 21786
rect 28974 21734 28986 21786
rect 29038 21734 29050 21786
rect 29102 21734 29114 21786
rect 29166 21734 29178 21786
rect 29230 21734 29242 21786
rect 29294 21734 31832 21786
rect 1104 21712 31832 21734
rect 5350 21632 5356 21684
rect 5408 21632 5414 21684
rect 6546 21632 6552 21684
rect 6604 21672 6610 21684
rect 6733 21675 6791 21681
rect 6733 21672 6745 21675
rect 6604 21644 6745 21672
rect 6604 21632 6610 21644
rect 6733 21641 6745 21644
rect 6779 21641 6791 21675
rect 6733 21635 6791 21641
rect 6825 21675 6883 21681
rect 6825 21641 6837 21675
rect 6871 21672 6883 21675
rect 7098 21672 7104 21684
rect 6871 21644 7104 21672
rect 6871 21641 6883 21644
rect 6825 21635 6883 21641
rect 5368 21604 5396 21632
rect 4816 21576 5396 21604
rect 4816 21545 4844 21576
rect 5534 21564 5540 21616
rect 5592 21604 5598 21616
rect 6086 21604 6092 21616
rect 5592 21576 6092 21604
rect 5592 21564 5598 21576
rect 6086 21564 6092 21576
rect 6144 21604 6150 21616
rect 6840 21604 6868 21635
rect 7098 21632 7104 21644
rect 7156 21672 7162 21684
rect 7156 21644 9444 21672
rect 7156 21632 7162 21644
rect 6144 21576 6868 21604
rect 6144 21564 6150 21576
rect 8662 21564 8668 21616
rect 8720 21564 8726 21616
rect 8754 21564 8760 21616
rect 8812 21604 8818 21616
rect 9309 21607 9367 21613
rect 9309 21604 9321 21607
rect 8812 21576 9321 21604
rect 8812 21564 8818 21576
rect 9309 21573 9321 21576
rect 9355 21573 9367 21607
rect 9416 21604 9444 21644
rect 9582 21632 9588 21684
rect 9640 21632 9646 21684
rect 10778 21632 10784 21684
rect 10836 21672 10842 21684
rect 11333 21675 11391 21681
rect 11333 21672 11345 21675
rect 10836 21644 11345 21672
rect 10836 21632 10842 21644
rect 11333 21641 11345 21644
rect 11379 21641 11391 21675
rect 11333 21635 11391 21641
rect 10220 21607 10278 21613
rect 9416 21576 10185 21604
rect 9309 21567 9367 21573
rect 4801 21539 4859 21545
rect 4801 21505 4813 21539
rect 4847 21505 4859 21539
rect 4801 21499 4859 21505
rect 5068 21539 5126 21545
rect 5068 21505 5080 21539
rect 5114 21536 5126 21539
rect 6178 21536 6184 21548
rect 5114 21508 6184 21536
rect 5114 21505 5126 21508
rect 5068 21499 5126 21505
rect 6178 21496 6184 21508
rect 6236 21496 6242 21548
rect 7374 21536 7380 21548
rect 7024 21508 7380 21536
rect 7024 21477 7052 21508
rect 7374 21496 7380 21508
rect 7432 21536 7438 21548
rect 7834 21536 7840 21548
rect 7432 21508 7840 21536
rect 7432 21496 7438 21508
rect 7834 21496 7840 21508
rect 7892 21496 7898 21548
rect 7929 21539 7987 21545
rect 7929 21505 7941 21539
rect 7975 21536 7987 21539
rect 8202 21536 8208 21548
rect 7975 21508 8208 21536
rect 7975 21505 7987 21508
rect 7929 21499 7987 21505
rect 8202 21496 8208 21508
rect 8260 21496 8266 21548
rect 8846 21496 8852 21548
rect 8904 21536 8910 21548
rect 9490 21545 9496 21548
rect 8941 21539 8999 21545
rect 8941 21536 8953 21539
rect 8904 21508 8953 21536
rect 8904 21496 8910 21508
rect 8941 21505 8953 21508
rect 8987 21505 8999 21539
rect 8941 21499 8999 21505
rect 9034 21539 9092 21545
rect 9034 21505 9046 21539
rect 9080 21505 9092 21539
rect 9034 21499 9092 21505
rect 9217 21539 9275 21545
rect 9217 21505 9229 21539
rect 9263 21536 9275 21539
rect 9447 21539 9496 21545
rect 9263 21508 9352 21536
rect 9263 21505 9275 21508
rect 9217 21499 9275 21505
rect 7009 21471 7067 21477
rect 7009 21437 7021 21471
rect 7055 21437 7067 21471
rect 7009 21431 7067 21437
rect 7190 21428 7196 21480
rect 7248 21468 7254 21480
rect 9048 21468 9076 21499
rect 7248 21440 9076 21468
rect 9324 21468 9352 21508
rect 9447 21505 9459 21539
rect 9493 21505 9496 21539
rect 9447 21499 9496 21505
rect 9490 21496 9496 21499
rect 9548 21496 9554 21548
rect 9953 21539 10011 21545
rect 9953 21505 9965 21539
rect 9999 21536 10011 21539
rect 10042 21536 10048 21548
rect 9999 21508 10048 21536
rect 9999 21505 10011 21508
rect 9953 21499 10011 21505
rect 10042 21496 10048 21508
rect 10100 21496 10106 21548
rect 10157 21536 10185 21576
rect 10220 21573 10232 21607
rect 10266 21604 10278 21607
rect 10410 21604 10416 21616
rect 10266 21576 10416 21604
rect 10266 21573 10278 21576
rect 10220 21567 10278 21573
rect 10410 21564 10416 21576
rect 10468 21564 10474 21616
rect 11348 21536 11376 21635
rect 12710 21632 12716 21684
rect 12768 21632 12774 21684
rect 13173 21675 13231 21681
rect 13173 21641 13185 21675
rect 13219 21672 13231 21675
rect 17497 21675 17555 21681
rect 13219 21644 13492 21672
rect 13219 21641 13231 21644
rect 13173 21635 13231 21641
rect 12069 21539 12127 21545
rect 12069 21536 12081 21539
rect 10157 21508 11008 21536
rect 11348 21508 12081 21536
rect 9858 21468 9864 21480
rect 9324 21440 9864 21468
rect 7248 21428 7254 21440
rect 6181 21403 6239 21409
rect 6181 21369 6193 21403
rect 6227 21400 6239 21403
rect 7208 21400 7236 21428
rect 6227 21372 7236 21400
rect 6227 21369 6239 21372
rect 6181 21363 6239 21369
rect 9324 21344 9352 21440
rect 9858 21428 9864 21440
rect 9916 21428 9922 21480
rect 10980 21468 11008 21508
rect 12069 21505 12081 21508
rect 12115 21505 12127 21539
rect 12805 21539 12863 21545
rect 12069 21499 12127 21505
rect 12176 21508 12756 21536
rect 12176 21468 12204 21508
rect 10980 21440 12204 21468
rect 12529 21471 12587 21477
rect 12529 21437 12541 21471
rect 12575 21468 12587 21471
rect 12728 21468 12756 21508
rect 12805 21505 12817 21539
rect 12851 21536 12863 21539
rect 13354 21536 13360 21548
rect 12851 21508 13360 21536
rect 12851 21505 12863 21508
rect 12805 21499 12863 21505
rect 13354 21496 13360 21508
rect 13412 21496 13418 21548
rect 13464 21545 13492 21644
rect 17497 21641 17509 21675
rect 17543 21672 17555 21675
rect 17586 21672 17592 21684
rect 17543 21644 17592 21672
rect 17543 21641 17555 21644
rect 17497 21635 17555 21641
rect 17586 21632 17592 21644
rect 17644 21632 17650 21684
rect 23474 21632 23480 21684
rect 23532 21632 23538 21684
rect 24489 21675 24547 21681
rect 24489 21641 24501 21675
rect 24535 21672 24547 21675
rect 24535 21644 24716 21672
rect 24535 21641 24547 21644
rect 24489 21635 24547 21641
rect 23842 21604 23848 21616
rect 19306 21576 23848 21604
rect 13449 21539 13507 21545
rect 13449 21505 13461 21539
rect 13495 21505 13507 21539
rect 13449 21499 13507 21505
rect 17589 21539 17647 21545
rect 17589 21505 17601 21539
rect 17635 21536 17647 21539
rect 18598 21536 18604 21548
rect 17635 21508 18604 21536
rect 17635 21505 17647 21508
rect 17589 21499 17647 21505
rect 18598 21496 18604 21508
rect 18656 21496 18662 21548
rect 19306 21468 19334 21576
rect 23842 21564 23848 21576
rect 23900 21564 23906 21616
rect 24118 21564 24124 21616
rect 24176 21564 24182 21616
rect 24210 21564 24216 21616
rect 24268 21604 24274 21616
rect 24268 21576 24624 21604
rect 24268 21564 24274 21576
rect 23658 21496 23664 21548
rect 23716 21496 23722 21548
rect 23937 21539 23995 21545
rect 23937 21505 23949 21539
rect 23983 21505 23995 21539
rect 23937 21499 23995 21505
rect 12575 21440 12609 21468
rect 12728 21440 19334 21468
rect 23952 21468 23980 21499
rect 24302 21496 24308 21548
rect 24360 21496 24366 21548
rect 24596 21545 24624 21576
rect 24581 21539 24639 21545
rect 24581 21505 24593 21539
rect 24627 21505 24639 21539
rect 24688 21536 24716 21644
rect 24762 21632 24768 21684
rect 24820 21672 24826 21684
rect 25225 21675 25283 21681
rect 25225 21672 25237 21675
rect 24820 21644 25237 21672
rect 24820 21632 24826 21644
rect 25225 21641 25237 21644
rect 25271 21641 25283 21675
rect 25225 21635 25283 21641
rect 29546 21632 29552 21684
rect 29604 21632 29610 21684
rect 24854 21564 24860 21616
rect 24912 21604 24918 21616
rect 25314 21604 25320 21616
rect 24912 21576 25320 21604
rect 24912 21564 24918 21576
rect 25314 21564 25320 21576
rect 25372 21564 25378 21616
rect 26050 21564 26056 21616
rect 26108 21564 26114 21616
rect 27430 21564 27436 21616
rect 27488 21604 27494 21616
rect 29457 21607 29515 21613
rect 29457 21604 29469 21607
rect 27488 21576 29469 21604
rect 27488 21564 27494 21576
rect 29457 21573 29469 21576
rect 29503 21573 29515 21607
rect 29457 21567 29515 21573
rect 26973 21539 27031 21545
rect 26973 21536 26985 21539
rect 24688 21508 26985 21536
rect 24581 21499 24639 21505
rect 26973 21505 26985 21508
rect 27019 21505 27031 21539
rect 26973 21499 27031 21505
rect 27249 21539 27307 21545
rect 27249 21505 27261 21539
rect 27295 21536 27307 21539
rect 27982 21536 27988 21548
rect 27295 21508 27988 21536
rect 27295 21505 27307 21508
rect 27249 21499 27307 21505
rect 27982 21496 27988 21508
rect 28040 21496 28046 21548
rect 30929 21539 30987 21545
rect 30929 21536 30941 21539
rect 29932 21508 30941 21536
rect 24670 21468 24676 21480
rect 23952 21440 24676 21468
rect 12575 21437 12587 21440
rect 12529 21431 12587 21437
rect 12544 21400 12572 21431
rect 24670 21428 24676 21440
rect 24728 21428 24734 21480
rect 26786 21428 26792 21480
rect 26844 21468 26850 21480
rect 27065 21471 27123 21477
rect 27065 21468 27077 21471
rect 26844 21440 27077 21468
rect 26844 21428 26850 21440
rect 27065 21437 27077 21440
rect 27111 21437 27123 21471
rect 27065 21431 27123 21437
rect 29365 21471 29423 21477
rect 29365 21437 29377 21471
rect 29411 21468 29423 21471
rect 29822 21468 29828 21480
rect 29411 21440 29828 21468
rect 29411 21437 29423 21440
rect 29365 21431 29423 21437
rect 29822 21428 29828 21440
rect 29880 21428 29886 21480
rect 12802 21400 12808 21412
rect 10980 21372 12808 21400
rect 6362 21292 6368 21344
rect 6420 21292 6426 21344
rect 9306 21292 9312 21344
rect 9364 21292 9370 21344
rect 10686 21292 10692 21344
rect 10744 21332 10750 21344
rect 10980 21332 11008 21372
rect 12802 21360 12808 21372
rect 12860 21360 12866 21412
rect 29932 21409 29960 21508
rect 30929 21505 30941 21508
rect 30975 21505 30987 21539
rect 30929 21499 30987 21505
rect 30098 21428 30104 21480
rect 30156 21468 30162 21480
rect 30561 21471 30619 21477
rect 30561 21468 30573 21471
rect 30156 21440 30573 21468
rect 30156 21428 30162 21440
rect 30561 21437 30573 21440
rect 30607 21437 30619 21471
rect 30561 21431 30619 21437
rect 29917 21403 29975 21409
rect 19306 21372 27476 21400
rect 10744 21304 11008 21332
rect 10744 21292 10750 21304
rect 11514 21292 11520 21344
rect 11572 21292 11578 21344
rect 13262 21292 13268 21344
rect 13320 21292 13326 21344
rect 17310 21292 17316 21344
rect 17368 21332 17374 21344
rect 19306 21332 19334 21372
rect 17368 21304 19334 21332
rect 17368 21292 17374 21304
rect 26970 21292 26976 21344
rect 27028 21292 27034 21344
rect 27448 21341 27476 21372
rect 29917 21369 29929 21403
rect 29963 21369 29975 21403
rect 29917 21363 29975 21369
rect 27433 21335 27491 21341
rect 27433 21301 27445 21335
rect 27479 21301 27491 21335
rect 27433 21295 27491 21301
rect 28994 21292 29000 21344
rect 29052 21332 29058 21344
rect 30009 21335 30067 21341
rect 30009 21332 30021 21335
rect 29052 21304 30021 21332
rect 29052 21292 29058 21304
rect 30009 21301 30021 21304
rect 30055 21301 30067 21335
rect 30009 21295 30067 21301
rect 30650 21292 30656 21344
rect 30708 21332 30714 21344
rect 30745 21335 30803 21341
rect 30745 21332 30757 21335
rect 30708 21304 30757 21332
rect 30708 21292 30714 21304
rect 30745 21301 30757 21304
rect 30791 21301 30803 21335
rect 30745 21295 30803 21301
rect 1104 21242 31832 21264
rect 1104 21190 4182 21242
rect 4234 21190 4246 21242
rect 4298 21190 4310 21242
rect 4362 21190 4374 21242
rect 4426 21190 4438 21242
rect 4490 21190 4502 21242
rect 4554 21190 10182 21242
rect 10234 21190 10246 21242
rect 10298 21190 10310 21242
rect 10362 21190 10374 21242
rect 10426 21190 10438 21242
rect 10490 21190 10502 21242
rect 10554 21190 16182 21242
rect 16234 21190 16246 21242
rect 16298 21190 16310 21242
rect 16362 21190 16374 21242
rect 16426 21190 16438 21242
rect 16490 21190 16502 21242
rect 16554 21190 22182 21242
rect 22234 21190 22246 21242
rect 22298 21190 22310 21242
rect 22362 21190 22374 21242
rect 22426 21190 22438 21242
rect 22490 21190 22502 21242
rect 22554 21190 28182 21242
rect 28234 21190 28246 21242
rect 28298 21190 28310 21242
rect 28362 21190 28374 21242
rect 28426 21190 28438 21242
rect 28490 21190 28502 21242
rect 28554 21190 31832 21242
rect 1104 21168 31832 21190
rect 5445 21131 5503 21137
rect 5445 21097 5457 21131
rect 5491 21128 5503 21131
rect 5626 21128 5632 21140
rect 5491 21100 5632 21128
rect 5491 21097 5503 21100
rect 5445 21091 5503 21097
rect 5626 21088 5632 21100
rect 5684 21088 5690 21140
rect 6178 21088 6184 21140
rect 6236 21088 6242 21140
rect 6362 21088 6368 21140
rect 6420 21088 6426 21140
rect 8938 21088 8944 21140
rect 8996 21088 9002 21140
rect 10594 21088 10600 21140
rect 10652 21088 10658 21140
rect 12526 21088 12532 21140
rect 12584 21128 12590 21140
rect 15286 21128 15292 21140
rect 12584 21100 15292 21128
rect 12584 21088 12590 21100
rect 15286 21088 15292 21100
rect 15344 21088 15350 21140
rect 23842 21088 23848 21140
rect 23900 21088 23906 21140
rect 26605 21131 26663 21137
rect 26605 21097 26617 21131
rect 26651 21128 26663 21131
rect 26970 21128 26976 21140
rect 26651 21100 26976 21128
rect 26651 21097 26663 21100
rect 26605 21091 26663 21097
rect 26970 21088 26976 21100
rect 27028 21088 27034 21140
rect 28261 21131 28319 21137
rect 28261 21097 28273 21131
rect 28307 21097 28319 21131
rect 28261 21091 28319 21097
rect 29549 21131 29607 21137
rect 29549 21097 29561 21131
rect 29595 21128 29607 21131
rect 29638 21128 29644 21140
rect 29595 21100 29644 21128
rect 29595 21097 29607 21100
rect 29549 21091 29607 21097
rect 6089 20995 6147 21001
rect 6089 20961 6101 20995
rect 6135 20992 6147 20995
rect 6270 20992 6276 21004
rect 6135 20964 6276 20992
rect 6135 20961 6147 20964
rect 6089 20955 6147 20961
rect 6270 20952 6276 20964
rect 6328 20952 6334 21004
rect 6380 20933 6408 21088
rect 10042 21020 10048 21072
rect 10100 21060 10106 21072
rect 10962 21060 10968 21072
rect 10100 21032 10968 21060
rect 10100 21020 10106 21032
rect 10962 21020 10968 21032
rect 11020 21020 11026 21072
rect 11514 21060 11520 21072
rect 11072 21032 11520 21060
rect 9585 20995 9643 21001
rect 9585 20961 9597 20995
rect 9631 20992 9643 20995
rect 9674 20992 9680 21004
rect 9631 20964 9680 20992
rect 9631 20961 9643 20964
rect 9585 20955 9643 20961
rect 9674 20952 9680 20964
rect 9732 20992 9738 21004
rect 10870 20992 10876 21004
rect 9732 20964 10876 20992
rect 9732 20952 9738 20964
rect 10870 20952 10876 20964
rect 10928 20952 10934 21004
rect 6365 20927 6423 20933
rect 6365 20893 6377 20927
rect 6411 20893 6423 20927
rect 6365 20887 6423 20893
rect 8478 20884 8484 20936
rect 8536 20933 8542 20936
rect 8536 20887 8548 20933
rect 8757 20927 8815 20933
rect 8757 20893 8769 20927
rect 8803 20924 8815 20927
rect 9858 20924 9864 20936
rect 8803 20896 9864 20924
rect 8803 20893 8815 20896
rect 8757 20887 8815 20893
rect 8536 20884 8542 20887
rect 9858 20884 9864 20896
rect 9916 20884 9922 20936
rect 10965 20927 11023 20933
rect 10965 20893 10977 20927
rect 11011 20924 11023 20927
rect 11072 20924 11100 21032
rect 11514 21020 11520 21032
rect 11572 21020 11578 21072
rect 23860 21060 23888 21088
rect 28074 21060 28080 21072
rect 23860 21032 28080 21060
rect 28074 21020 28080 21032
rect 28132 21020 28138 21072
rect 11149 20995 11207 21001
rect 11149 20961 11161 20995
rect 11195 20992 11207 20995
rect 11422 20992 11428 21004
rect 11195 20964 11428 20992
rect 11195 20961 11207 20964
rect 11149 20955 11207 20961
rect 11422 20952 11428 20964
rect 11480 20992 11486 21004
rect 12250 20992 12256 21004
rect 11480 20964 12256 20992
rect 11480 20952 11486 20964
rect 12250 20952 12256 20964
rect 12308 20992 12314 21004
rect 14918 20992 14924 21004
rect 12308 20964 14924 20992
rect 12308 20952 12314 20964
rect 14918 20952 14924 20964
rect 14976 20952 14982 21004
rect 24946 20952 24952 21004
rect 25004 20992 25010 21004
rect 25004 20964 27016 20992
rect 25004 20952 25010 20964
rect 11011 20896 11100 20924
rect 11011 20893 11023 20896
rect 10965 20887 11023 20893
rect 11238 20884 11244 20936
rect 11296 20884 11302 20936
rect 11330 20884 11336 20936
rect 11388 20924 11394 20936
rect 12158 20924 12164 20936
rect 11388 20896 12164 20924
rect 11388 20884 11394 20896
rect 12158 20884 12164 20896
rect 12216 20884 12222 20936
rect 14182 20924 14188 20936
rect 12406 20896 14188 20924
rect 8386 20816 8392 20868
rect 8444 20856 8450 20868
rect 9214 20856 9220 20868
rect 8444 20828 9220 20856
rect 8444 20816 8450 20828
rect 9214 20816 9220 20828
rect 9272 20856 9278 20868
rect 9401 20859 9459 20865
rect 9401 20856 9413 20859
rect 9272 20828 9413 20856
rect 9272 20816 9278 20828
rect 9401 20825 9413 20828
rect 9447 20856 9459 20859
rect 11057 20859 11115 20865
rect 11057 20856 11069 20859
rect 9447 20828 11069 20856
rect 9447 20825 9459 20828
rect 9401 20819 9459 20825
rect 11057 20825 11069 20828
rect 11103 20825 11115 20859
rect 11256 20856 11284 20884
rect 12406 20856 12434 20896
rect 14182 20884 14188 20896
rect 14240 20924 14246 20936
rect 14277 20927 14335 20933
rect 14277 20924 14289 20927
rect 14240 20896 14289 20924
rect 14240 20884 14246 20896
rect 14277 20893 14289 20896
rect 14323 20893 14335 20927
rect 14277 20887 14335 20893
rect 25038 20884 25044 20936
rect 25096 20924 25102 20936
rect 25869 20927 25927 20933
rect 25869 20924 25881 20927
rect 25096 20896 25881 20924
rect 25096 20884 25102 20896
rect 25869 20893 25881 20896
rect 25915 20924 25927 20927
rect 26053 20927 26111 20933
rect 26053 20924 26065 20927
rect 25915 20896 26065 20924
rect 25915 20893 25927 20896
rect 25869 20887 25927 20893
rect 26053 20893 26065 20896
rect 26099 20893 26111 20927
rect 26053 20887 26111 20893
rect 26421 20927 26479 20933
rect 26421 20893 26433 20927
rect 26467 20924 26479 20927
rect 26510 20924 26516 20936
rect 26467 20896 26516 20924
rect 26467 20893 26479 20896
rect 26421 20887 26479 20893
rect 26510 20884 26516 20896
rect 26568 20884 26574 20936
rect 26988 20924 27016 20964
rect 27062 20952 27068 21004
rect 27120 20992 27126 21004
rect 27525 20995 27583 21001
rect 27525 20992 27537 20995
rect 27120 20964 27537 20992
rect 27120 20952 27126 20964
rect 27525 20961 27537 20964
rect 27571 20961 27583 20995
rect 27525 20955 27583 20961
rect 27430 20924 27436 20936
rect 26988 20896 27436 20924
rect 27430 20884 27436 20896
rect 27488 20924 27494 20936
rect 28276 20924 28304 21091
rect 29638 21088 29644 21100
rect 29696 21088 29702 21140
rect 29748 21100 31248 21128
rect 29365 21063 29423 21069
rect 29365 21029 29377 21063
rect 29411 21060 29423 21063
rect 29748 21060 29776 21100
rect 29411 21032 29776 21060
rect 29411 21029 29423 21032
rect 29365 21023 29423 21029
rect 28813 20995 28871 21001
rect 28813 20961 28825 20995
rect 28859 20992 28871 20995
rect 29546 20992 29552 21004
rect 28859 20964 29552 20992
rect 28859 20961 28871 20964
rect 28813 20955 28871 20961
rect 29546 20952 29552 20964
rect 29604 20992 29610 21004
rect 29730 20992 29736 21004
rect 29604 20964 29736 20992
rect 29604 20952 29610 20964
rect 29730 20952 29736 20964
rect 29788 20952 29794 21004
rect 30852 20964 31156 20992
rect 28905 20927 28963 20933
rect 28905 20924 28917 20927
rect 27488 20896 28917 20924
rect 27488 20884 27494 20896
rect 28905 20893 28917 20896
rect 28951 20893 28963 20927
rect 28905 20887 28963 20893
rect 28994 20884 29000 20936
rect 29052 20884 29058 20936
rect 30650 20884 30656 20936
rect 30708 20933 30714 20936
rect 30708 20924 30720 20933
rect 30708 20896 30753 20924
rect 30708 20887 30720 20896
rect 30708 20884 30714 20887
rect 11256 20828 12434 20856
rect 11057 20819 11115 20825
rect 12894 20816 12900 20868
rect 12952 20816 12958 20868
rect 26237 20859 26295 20865
rect 26237 20825 26249 20859
rect 26283 20825 26295 20859
rect 26237 20819 26295 20825
rect 26329 20859 26387 20865
rect 26329 20825 26341 20859
rect 26375 20856 26387 20859
rect 27246 20856 27252 20868
rect 26375 20828 27252 20856
rect 26375 20825 26387 20828
rect 26329 20819 26387 20825
rect 7377 20791 7435 20797
rect 7377 20757 7389 20791
rect 7423 20788 7435 20791
rect 8754 20788 8760 20800
rect 7423 20760 8760 20788
rect 7423 20757 7435 20760
rect 7377 20751 7435 20757
rect 8754 20748 8760 20760
rect 8812 20748 8818 20800
rect 9306 20748 9312 20800
rect 9364 20748 9370 20800
rect 10870 20748 10876 20800
rect 10928 20788 10934 20800
rect 12618 20788 12624 20800
rect 10928 20760 12624 20788
rect 10928 20748 10934 20760
rect 12618 20748 12624 20760
rect 12676 20748 12682 20800
rect 14182 20748 14188 20800
rect 14240 20748 14246 20800
rect 25314 20748 25320 20800
rect 25372 20748 25378 20800
rect 26252 20788 26280 20819
rect 27246 20816 27252 20828
rect 27304 20816 27310 20868
rect 27341 20859 27399 20865
rect 27341 20825 27353 20859
rect 27387 20856 27399 20859
rect 27890 20856 27896 20868
rect 27387 20828 27896 20856
rect 27387 20825 27399 20828
rect 27341 20819 27399 20825
rect 27890 20816 27896 20828
rect 27948 20816 27954 20868
rect 28074 20816 28080 20868
rect 28132 20856 28138 20868
rect 28169 20859 28227 20865
rect 28169 20856 28181 20859
rect 28132 20828 28181 20856
rect 28132 20816 28138 20828
rect 28169 20825 28181 20828
rect 28215 20856 28227 20859
rect 28626 20856 28632 20868
rect 28215 20828 28632 20856
rect 28215 20825 28227 20828
rect 28169 20819 28227 20825
rect 28626 20816 28632 20828
rect 28684 20856 28690 20868
rect 30852 20856 30880 20964
rect 30929 20927 30987 20933
rect 30929 20893 30941 20927
rect 30975 20893 30987 20927
rect 30929 20887 30987 20893
rect 28684 20828 30880 20856
rect 28684 20816 28690 20828
rect 26694 20788 26700 20800
rect 26252 20760 26700 20788
rect 26694 20748 26700 20760
rect 26752 20748 26758 20800
rect 26970 20748 26976 20800
rect 27028 20748 27034 20800
rect 30558 20748 30564 20800
rect 30616 20788 30622 20800
rect 30944 20788 30972 20887
rect 31128 20868 31156 20964
rect 31220 20933 31248 21100
rect 31205 20927 31263 20933
rect 31205 20893 31217 20927
rect 31251 20893 31263 20927
rect 31205 20887 31263 20893
rect 31110 20816 31116 20868
rect 31168 20816 31174 20868
rect 30616 20760 30972 20788
rect 30616 20748 30622 20760
rect 31018 20748 31024 20800
rect 31076 20748 31082 20800
rect 1104 20698 31832 20720
rect 1104 20646 4922 20698
rect 4974 20646 4986 20698
rect 5038 20646 5050 20698
rect 5102 20646 5114 20698
rect 5166 20646 5178 20698
rect 5230 20646 5242 20698
rect 5294 20646 10922 20698
rect 10974 20646 10986 20698
rect 11038 20646 11050 20698
rect 11102 20646 11114 20698
rect 11166 20646 11178 20698
rect 11230 20646 11242 20698
rect 11294 20646 16922 20698
rect 16974 20646 16986 20698
rect 17038 20646 17050 20698
rect 17102 20646 17114 20698
rect 17166 20646 17178 20698
rect 17230 20646 17242 20698
rect 17294 20646 22922 20698
rect 22974 20646 22986 20698
rect 23038 20646 23050 20698
rect 23102 20646 23114 20698
rect 23166 20646 23178 20698
rect 23230 20646 23242 20698
rect 23294 20646 28922 20698
rect 28974 20646 28986 20698
rect 29038 20646 29050 20698
rect 29102 20646 29114 20698
rect 29166 20646 29178 20698
rect 29230 20646 29242 20698
rect 29294 20646 31832 20698
rect 1104 20624 31832 20646
rect 9217 20587 9275 20593
rect 9217 20553 9229 20587
rect 9263 20584 9275 20587
rect 9306 20584 9312 20596
rect 9263 20556 9312 20584
rect 9263 20553 9275 20556
rect 9217 20547 9275 20553
rect 9306 20544 9312 20556
rect 9364 20544 9370 20596
rect 10778 20544 10784 20596
rect 10836 20584 10842 20596
rect 11422 20584 11428 20596
rect 10836 20556 11428 20584
rect 10836 20544 10842 20556
rect 11422 20544 11428 20556
rect 11480 20544 11486 20596
rect 13354 20544 13360 20596
rect 13412 20584 13418 20596
rect 14645 20587 14703 20593
rect 14645 20584 14657 20587
rect 13412 20556 14657 20584
rect 13412 20544 13418 20556
rect 14645 20553 14657 20556
rect 14691 20584 14703 20587
rect 14691 20556 22094 20584
rect 14691 20553 14703 20556
rect 14645 20547 14703 20553
rect 8294 20476 8300 20528
rect 8352 20516 8358 20528
rect 8481 20519 8539 20525
rect 8481 20516 8493 20519
rect 8352 20488 8493 20516
rect 8352 20476 8358 20488
rect 8481 20485 8493 20488
rect 8527 20485 8539 20519
rect 13173 20519 13231 20525
rect 8481 20479 8539 20485
rect 8588 20488 9904 20516
rect 7466 20408 7472 20460
rect 7524 20408 7530 20460
rect 7742 20408 7748 20460
rect 7800 20448 7806 20460
rect 8588 20448 8616 20488
rect 7800 20420 8616 20448
rect 8665 20451 8723 20457
rect 7800 20408 7806 20420
rect 8665 20417 8677 20451
rect 8711 20448 8723 20451
rect 8754 20448 8760 20460
rect 8711 20420 8760 20448
rect 8711 20417 8723 20420
rect 8665 20411 8723 20417
rect 8754 20408 8760 20420
rect 8812 20408 8818 20460
rect 9490 20408 9496 20460
rect 9548 20408 9554 20460
rect 9585 20451 9643 20457
rect 9585 20417 9597 20451
rect 9631 20417 9643 20451
rect 9585 20411 9643 20417
rect 9677 20451 9735 20457
rect 9677 20417 9689 20451
rect 9723 20448 9735 20451
rect 9766 20448 9772 20460
rect 9723 20420 9772 20448
rect 9723 20417 9735 20420
rect 9677 20411 9735 20417
rect 6914 20340 6920 20392
rect 6972 20380 6978 20392
rect 7653 20383 7711 20389
rect 7653 20380 7665 20383
rect 6972 20352 7665 20380
rect 6972 20340 6978 20352
rect 7653 20349 7665 20352
rect 7699 20349 7711 20383
rect 7653 20343 7711 20349
rect 8846 20340 8852 20392
rect 8904 20340 8910 20392
rect 9600 20380 9628 20411
rect 9508 20352 9628 20380
rect 8864 20312 8892 20340
rect 9309 20315 9367 20321
rect 9309 20312 9321 20315
rect 8864 20284 9321 20312
rect 9309 20281 9321 20284
rect 9355 20281 9367 20315
rect 9309 20275 9367 20281
rect 9508 20256 9536 20352
rect 7282 20204 7288 20256
rect 7340 20204 7346 20256
rect 9490 20204 9496 20256
rect 9548 20204 9554 20256
rect 9692 20244 9720 20411
rect 9766 20408 9772 20420
rect 9824 20408 9830 20460
rect 9876 20457 9904 20488
rect 13173 20485 13185 20519
rect 13219 20516 13231 20519
rect 13262 20516 13268 20528
rect 13219 20488 13268 20516
rect 13219 20485 13231 20488
rect 13173 20479 13231 20485
rect 13262 20476 13268 20488
rect 13320 20476 13326 20528
rect 14182 20476 14188 20528
rect 14240 20476 14246 20528
rect 9861 20451 9919 20457
rect 9861 20417 9873 20451
rect 9907 20417 9919 20451
rect 9861 20411 9919 20417
rect 11514 20340 11520 20392
rect 11572 20380 11578 20392
rect 12894 20380 12900 20392
rect 11572 20352 12900 20380
rect 11572 20340 11578 20352
rect 12894 20340 12900 20352
rect 12952 20340 12958 20392
rect 9766 20272 9772 20324
rect 9824 20312 9830 20324
rect 12526 20312 12532 20324
rect 9824 20284 12532 20312
rect 9824 20272 9830 20284
rect 12526 20272 12532 20284
rect 12584 20272 12590 20324
rect 12342 20244 12348 20256
rect 9692 20216 12348 20244
rect 12342 20204 12348 20216
rect 12400 20204 12406 20256
rect 12912 20244 12940 20340
rect 14550 20244 14556 20256
rect 12912 20216 14556 20244
rect 14550 20204 14556 20216
rect 14608 20204 14614 20256
rect 22066 20244 22094 20556
rect 25038 20544 25044 20596
rect 25096 20544 25102 20596
rect 25314 20544 25320 20596
rect 25372 20584 25378 20596
rect 25501 20587 25559 20593
rect 25501 20584 25513 20587
rect 25372 20556 25513 20584
rect 25372 20544 25378 20556
rect 25501 20553 25513 20556
rect 25547 20553 25559 20587
rect 25501 20547 25559 20553
rect 26970 20544 26976 20596
rect 27028 20544 27034 20596
rect 27890 20544 27896 20596
rect 27948 20544 27954 20596
rect 28994 20544 29000 20596
rect 29052 20584 29058 20596
rect 29273 20587 29331 20593
rect 29273 20584 29285 20587
rect 29052 20556 29285 20584
rect 29052 20544 29058 20556
rect 29273 20553 29285 20556
rect 29319 20584 29331 20587
rect 30098 20584 30104 20596
rect 29319 20556 30104 20584
rect 29319 20553 29331 20556
rect 29273 20547 29331 20553
rect 30098 20544 30104 20556
rect 30156 20544 30162 20596
rect 26142 20516 26148 20528
rect 23676 20488 26148 20516
rect 23676 20457 23704 20488
rect 26142 20476 26148 20488
rect 26200 20476 26206 20528
rect 23934 20457 23940 20460
rect 23661 20451 23719 20457
rect 23661 20417 23673 20451
rect 23707 20417 23719 20451
rect 23661 20411 23719 20417
rect 23928 20411 23940 20457
rect 23934 20408 23940 20411
rect 23992 20408 23998 20460
rect 24946 20408 24952 20460
rect 25004 20448 25010 20460
rect 25593 20451 25651 20457
rect 25593 20448 25605 20451
rect 25004 20420 25605 20448
rect 25004 20408 25010 20420
rect 25593 20417 25605 20420
rect 25639 20417 25651 20451
rect 25593 20411 25651 20417
rect 26513 20451 26571 20457
rect 26513 20417 26525 20451
rect 26559 20448 26571 20451
rect 26988 20448 27016 20544
rect 27246 20476 27252 20528
rect 27304 20476 27310 20528
rect 30408 20519 30466 20525
rect 30408 20485 30420 20519
rect 30454 20516 30466 20519
rect 31018 20516 31024 20528
rect 30454 20488 31024 20516
rect 30454 20485 30466 20488
rect 30408 20479 30466 20485
rect 31018 20476 31024 20488
rect 31076 20476 31082 20528
rect 26559 20420 27016 20448
rect 27264 20448 27292 20476
rect 28445 20451 28503 20457
rect 28445 20448 28457 20451
rect 27264 20420 28457 20448
rect 26559 20417 26571 20420
rect 26513 20411 26571 20417
rect 28445 20417 28457 20420
rect 28491 20417 28503 20451
rect 28445 20411 28503 20417
rect 30558 20408 30564 20460
rect 30616 20448 30622 20460
rect 30653 20451 30711 20457
rect 30653 20448 30665 20451
rect 30616 20420 30665 20448
rect 30616 20408 30622 20420
rect 30653 20417 30665 20420
rect 30699 20417 30711 20451
rect 30653 20411 30711 20417
rect 25222 20340 25228 20392
rect 25280 20380 25286 20392
rect 25685 20383 25743 20389
rect 25685 20380 25697 20383
rect 25280 20352 25697 20380
rect 25280 20340 25286 20352
rect 25685 20349 25697 20352
rect 25731 20349 25743 20383
rect 25685 20343 25743 20349
rect 26234 20340 26240 20392
rect 26292 20380 26298 20392
rect 26973 20383 27031 20389
rect 26973 20380 26985 20383
rect 26292 20352 26985 20380
rect 26292 20340 26298 20352
rect 26973 20349 26985 20352
rect 27019 20349 27031 20383
rect 26973 20343 27031 20349
rect 27249 20383 27307 20389
rect 27249 20349 27261 20383
rect 27295 20380 27307 20383
rect 27295 20352 29408 20380
rect 27295 20349 27307 20352
rect 27249 20343 27307 20349
rect 29380 20324 29408 20352
rect 24596 20284 26464 20312
rect 24596 20244 24624 20284
rect 22066 20216 24624 20244
rect 25130 20204 25136 20256
rect 25188 20204 25194 20256
rect 26326 20204 26332 20256
rect 26384 20204 26390 20256
rect 26436 20244 26464 20284
rect 29362 20272 29368 20324
rect 29420 20272 29426 20324
rect 31202 20244 31208 20256
rect 26436 20216 31208 20244
rect 31202 20204 31208 20216
rect 31260 20204 31266 20256
rect 1104 20154 31832 20176
rect 1104 20102 4182 20154
rect 4234 20102 4246 20154
rect 4298 20102 4310 20154
rect 4362 20102 4374 20154
rect 4426 20102 4438 20154
rect 4490 20102 4502 20154
rect 4554 20102 10182 20154
rect 10234 20102 10246 20154
rect 10298 20102 10310 20154
rect 10362 20102 10374 20154
rect 10426 20102 10438 20154
rect 10490 20102 10502 20154
rect 10554 20102 16182 20154
rect 16234 20102 16246 20154
rect 16298 20102 16310 20154
rect 16362 20102 16374 20154
rect 16426 20102 16438 20154
rect 16490 20102 16502 20154
rect 16554 20102 22182 20154
rect 22234 20102 22246 20154
rect 22298 20102 22310 20154
rect 22362 20102 22374 20154
rect 22426 20102 22438 20154
rect 22490 20102 22502 20154
rect 22554 20102 28182 20154
rect 28234 20102 28246 20154
rect 28298 20102 28310 20154
rect 28362 20102 28374 20154
rect 28426 20102 28438 20154
rect 28490 20102 28502 20154
rect 28554 20102 31832 20154
rect 1104 20080 31832 20102
rect 23934 20000 23940 20052
rect 23992 20040 23998 20052
rect 24029 20043 24087 20049
rect 24029 20040 24041 20043
rect 23992 20012 24041 20040
rect 23992 20000 23998 20012
rect 24029 20009 24041 20012
rect 24075 20009 24087 20043
rect 24029 20003 24087 20009
rect 25130 20000 25136 20052
rect 25188 20000 25194 20052
rect 27246 20000 27252 20052
rect 27304 20040 27310 20052
rect 27433 20043 27491 20049
rect 27433 20040 27445 20043
rect 27304 20012 27445 20040
rect 27304 20000 27310 20012
rect 27433 20009 27445 20012
rect 27479 20009 27491 20043
rect 27433 20003 27491 20009
rect 27982 20000 27988 20052
rect 28040 20040 28046 20052
rect 28537 20043 28595 20049
rect 28537 20040 28549 20043
rect 28040 20012 28549 20040
rect 28040 20000 28046 20012
rect 28537 20009 28549 20012
rect 28583 20009 28595 20043
rect 28537 20003 28595 20009
rect 31389 20043 31447 20049
rect 31389 20009 31401 20043
rect 31435 20040 31447 20043
rect 31435 20012 31892 20040
rect 31435 20009 31447 20012
rect 31389 20003 31447 20009
rect 8389 19975 8447 19981
rect 8389 19941 8401 19975
rect 8435 19941 8447 19975
rect 8389 19935 8447 19941
rect 4433 19907 4491 19913
rect 4433 19873 4445 19907
rect 4479 19904 4491 19907
rect 4706 19904 4712 19916
rect 4479 19876 4712 19904
rect 4479 19873 4491 19876
rect 4433 19867 4491 19873
rect 4706 19864 4712 19876
rect 4764 19904 4770 19916
rect 5810 19904 5816 19916
rect 4764 19876 5816 19904
rect 4764 19864 4770 19876
rect 5810 19864 5816 19876
rect 5868 19864 5874 19916
rect 8404 19904 8432 19935
rect 9490 19904 9496 19916
rect 8404 19876 9496 19904
rect 9490 19864 9496 19876
rect 9548 19864 9554 19916
rect 18966 19864 18972 19916
rect 19024 19904 19030 19916
rect 20438 19904 20444 19916
rect 19024 19876 20444 19904
rect 19024 19864 19030 19876
rect 20438 19864 20444 19876
rect 20496 19864 20502 19916
rect 22002 19864 22008 19916
rect 22060 19864 22066 19916
rect 5445 19839 5503 19845
rect 5445 19805 5457 19839
rect 5491 19836 5503 19839
rect 5534 19836 5540 19848
rect 5491 19808 5540 19836
rect 5491 19805 5503 19808
rect 5445 19799 5503 19805
rect 5534 19796 5540 19808
rect 5592 19796 5598 19848
rect 6914 19796 6920 19848
rect 6972 19836 6978 19848
rect 7282 19845 7288 19848
rect 7009 19839 7067 19845
rect 7009 19836 7021 19839
rect 6972 19808 7021 19836
rect 6972 19796 6978 19808
rect 7009 19805 7021 19808
rect 7055 19805 7067 19839
rect 7276 19836 7288 19845
rect 7243 19808 7288 19836
rect 7009 19799 7067 19805
rect 7276 19799 7288 19808
rect 7282 19796 7288 19799
rect 7340 19796 7346 19848
rect 11977 19839 12035 19845
rect 11977 19805 11989 19839
rect 12023 19836 12035 19839
rect 12158 19836 12164 19848
rect 12023 19808 12164 19836
rect 12023 19805 12035 19808
rect 11977 19799 12035 19805
rect 12158 19796 12164 19808
rect 12216 19796 12222 19848
rect 12250 19796 12256 19848
rect 12308 19796 12314 19848
rect 12894 19796 12900 19848
rect 12952 19836 12958 19848
rect 13357 19839 13415 19845
rect 13357 19836 13369 19839
rect 12952 19808 13369 19836
rect 12952 19796 12958 19808
rect 13357 19805 13369 19808
rect 13403 19805 13415 19839
rect 13357 19799 13415 19805
rect 17678 19796 17684 19848
rect 17736 19796 17742 19848
rect 20714 19796 20720 19848
rect 20772 19796 20778 19848
rect 21174 19796 21180 19848
rect 21232 19796 21238 19848
rect 22830 19796 22836 19848
rect 22888 19796 22894 19848
rect 24213 19839 24271 19845
rect 24213 19805 24225 19839
rect 24259 19836 24271 19839
rect 25148 19836 25176 20000
rect 31864 19984 31892 20012
rect 31846 19932 31852 19984
rect 31904 19932 31910 19984
rect 24259 19808 25176 19836
rect 26053 19839 26111 19845
rect 24259 19805 24271 19808
rect 24213 19799 24271 19805
rect 26053 19805 26065 19839
rect 26099 19836 26111 19839
rect 26142 19836 26148 19848
rect 26099 19808 26148 19836
rect 26099 19805 26111 19808
rect 26053 19799 26111 19805
rect 26142 19796 26148 19808
rect 26200 19796 26206 19848
rect 26326 19845 26332 19848
rect 26320 19836 26332 19845
rect 26287 19808 26332 19836
rect 26320 19799 26332 19808
rect 26326 19796 26332 19799
rect 26384 19796 26390 19848
rect 28718 19845 28724 19848
rect 28716 19836 28724 19845
rect 28679 19808 28724 19836
rect 28716 19799 28724 19808
rect 28718 19796 28724 19799
rect 28776 19796 28782 19848
rect 28813 19839 28871 19845
rect 28813 19805 28825 19839
rect 28859 19836 28871 19839
rect 28994 19836 29000 19848
rect 28859 19808 29000 19836
rect 28859 19805 28871 19808
rect 28813 19799 28871 19805
rect 28994 19796 29000 19808
rect 29052 19796 29058 19848
rect 29088 19839 29146 19845
rect 29088 19805 29100 19839
rect 29134 19805 29146 19839
rect 29088 19799 29146 19805
rect 29181 19839 29239 19845
rect 29181 19805 29193 19839
rect 29227 19836 29239 19839
rect 29362 19836 29368 19848
rect 29227 19808 29368 19836
rect 29227 19805 29239 19808
rect 29181 19799 29239 19805
rect 4157 19771 4215 19777
rect 4157 19737 4169 19771
rect 4203 19768 4215 19771
rect 4801 19771 4859 19777
rect 4801 19768 4813 19771
rect 4203 19740 4813 19768
rect 4203 19737 4215 19740
rect 4157 19731 4215 19737
rect 4801 19737 4813 19740
rect 4847 19737 4859 19771
rect 4801 19731 4859 19737
rect 21821 19771 21879 19777
rect 21821 19737 21833 19771
rect 21867 19768 21879 19771
rect 22281 19771 22339 19777
rect 22281 19768 22293 19771
rect 21867 19740 22293 19768
rect 21867 19737 21879 19740
rect 21821 19731 21879 19737
rect 22281 19737 22293 19740
rect 22327 19737 22339 19771
rect 22281 19731 22339 19737
rect 22738 19728 22744 19780
rect 22796 19768 22802 19780
rect 23658 19768 23664 19780
rect 22796 19740 23664 19768
rect 22796 19728 22802 19740
rect 23658 19728 23664 19740
rect 23716 19768 23722 19780
rect 27338 19768 27344 19780
rect 23716 19740 27344 19768
rect 23716 19728 23722 19740
rect 27338 19728 27344 19740
rect 27396 19768 27402 19780
rect 28902 19768 28908 19780
rect 27396 19740 28908 19768
rect 27396 19728 27402 19740
rect 28902 19728 28908 19740
rect 28960 19728 28966 19780
rect 29104 19768 29132 19799
rect 29362 19796 29368 19808
rect 29420 19796 29426 19848
rect 29638 19796 29644 19848
rect 29696 19796 29702 19848
rect 31202 19796 31208 19848
rect 31260 19796 31266 19848
rect 29656 19768 29684 19796
rect 29104 19740 29684 19768
rect 3142 19660 3148 19712
rect 3200 19700 3206 19712
rect 3789 19703 3847 19709
rect 3789 19700 3801 19703
rect 3200 19672 3801 19700
rect 3200 19660 3206 19672
rect 3789 19669 3801 19672
rect 3835 19669 3847 19703
rect 3789 19663 3847 19669
rect 4249 19703 4307 19709
rect 4249 19669 4261 19703
rect 4295 19700 4307 19703
rect 4890 19700 4896 19712
rect 4295 19672 4896 19700
rect 4295 19669 4307 19672
rect 4249 19663 4307 19669
rect 4890 19660 4896 19672
rect 4948 19660 4954 19712
rect 8938 19660 8944 19712
rect 8996 19660 9002 19712
rect 11330 19660 11336 19712
rect 11388 19660 11394 19712
rect 12066 19660 12072 19712
rect 12124 19660 12130 19712
rect 12802 19660 12808 19712
rect 12860 19660 12866 19712
rect 17494 19660 17500 19712
rect 17552 19660 17558 19712
rect 18322 19660 18328 19712
rect 18380 19660 18386 19712
rect 20162 19660 20168 19712
rect 20220 19660 20226 19712
rect 20990 19660 20996 19712
rect 21048 19660 21054 19712
rect 21450 19660 21456 19712
rect 21508 19660 21514 19712
rect 21634 19660 21640 19712
rect 21692 19700 21698 19712
rect 21913 19703 21971 19709
rect 21913 19700 21925 19703
rect 21692 19672 21925 19700
rect 21692 19660 21698 19672
rect 21913 19669 21925 19672
rect 21959 19669 21971 19703
rect 28920 19700 28948 19728
rect 29454 19700 29460 19712
rect 28920 19672 29460 19700
rect 21913 19663 21971 19669
rect 29454 19660 29460 19672
rect 29512 19660 29518 19712
rect 1104 19610 31832 19632
rect 1104 19558 4922 19610
rect 4974 19558 4986 19610
rect 5038 19558 5050 19610
rect 5102 19558 5114 19610
rect 5166 19558 5178 19610
rect 5230 19558 5242 19610
rect 5294 19558 10922 19610
rect 10974 19558 10986 19610
rect 11038 19558 11050 19610
rect 11102 19558 11114 19610
rect 11166 19558 11178 19610
rect 11230 19558 11242 19610
rect 11294 19558 16922 19610
rect 16974 19558 16986 19610
rect 17038 19558 17050 19610
rect 17102 19558 17114 19610
rect 17166 19558 17178 19610
rect 17230 19558 17242 19610
rect 17294 19558 22922 19610
rect 22974 19558 22986 19610
rect 23038 19558 23050 19610
rect 23102 19558 23114 19610
rect 23166 19558 23178 19610
rect 23230 19558 23242 19610
rect 23294 19558 28922 19610
rect 28974 19558 28986 19610
rect 29038 19558 29050 19610
rect 29102 19558 29114 19610
rect 29166 19558 29178 19610
rect 29230 19558 29242 19610
rect 29294 19558 31832 19610
rect 1104 19536 31832 19558
rect 3881 19499 3939 19505
rect 3881 19465 3893 19499
rect 3927 19496 3939 19499
rect 5166 19496 5172 19508
rect 3927 19468 5172 19496
rect 3927 19465 3939 19468
rect 3881 19459 3939 19465
rect 5166 19456 5172 19468
rect 5224 19456 5230 19508
rect 5353 19499 5411 19505
rect 5353 19465 5365 19499
rect 5399 19496 5411 19499
rect 5534 19496 5540 19508
rect 5399 19468 5540 19496
rect 5399 19465 5411 19468
rect 5353 19459 5411 19465
rect 5534 19456 5540 19468
rect 5592 19456 5598 19508
rect 7466 19456 7472 19508
rect 7524 19496 7530 19508
rect 7837 19499 7895 19505
rect 7837 19496 7849 19499
rect 7524 19468 7849 19496
rect 7524 19456 7530 19468
rect 7837 19465 7849 19468
rect 7883 19465 7895 19499
rect 7837 19459 7895 19465
rect 8205 19499 8263 19505
rect 8205 19465 8217 19499
rect 8251 19496 8263 19499
rect 8938 19496 8944 19508
rect 8251 19468 8944 19496
rect 8251 19465 8263 19468
rect 8205 19459 8263 19465
rect 8938 19456 8944 19468
rect 8996 19456 9002 19508
rect 11333 19499 11391 19505
rect 11333 19465 11345 19499
rect 11379 19496 11391 19499
rect 11379 19468 11744 19496
rect 11379 19465 11391 19468
rect 11333 19459 11391 19465
rect 2516 19400 6960 19428
rect 2516 19369 2544 19400
rect 3988 19372 4016 19400
rect 2501 19363 2559 19369
rect 2501 19329 2513 19363
rect 2547 19329 2559 19363
rect 2501 19323 2559 19329
rect 2768 19363 2826 19369
rect 2768 19329 2780 19363
rect 2814 19360 2826 19363
rect 3050 19360 3056 19372
rect 2814 19332 3056 19360
rect 2814 19329 2826 19332
rect 2768 19323 2826 19329
rect 3050 19320 3056 19332
rect 3108 19320 3114 19372
rect 3970 19320 3976 19372
rect 4028 19320 4034 19372
rect 4246 19369 4252 19372
rect 4240 19323 4252 19369
rect 4246 19320 4252 19323
rect 4304 19320 4310 19372
rect 5994 19320 6000 19372
rect 6052 19320 6058 19372
rect 6380 19369 6408 19400
rect 6932 19372 6960 19400
rect 9968 19400 11560 19428
rect 6365 19363 6423 19369
rect 6365 19329 6377 19363
rect 6411 19329 6423 19363
rect 6621 19363 6679 19369
rect 6621 19360 6633 19363
rect 6365 19323 6423 19329
rect 6472 19332 6633 19360
rect 6472 19292 6500 19332
rect 6621 19329 6633 19332
rect 6667 19329 6679 19363
rect 6621 19323 6679 19329
rect 6914 19320 6920 19372
rect 6972 19320 6978 19372
rect 9858 19320 9864 19372
rect 9916 19360 9922 19372
rect 9968 19369 9996 19400
rect 11532 19372 11560 19400
rect 9953 19363 10011 19369
rect 9953 19360 9965 19363
rect 9916 19332 9965 19360
rect 9916 19320 9922 19332
rect 9953 19329 9965 19332
rect 9999 19329 10011 19363
rect 9953 19323 10011 19329
rect 10220 19363 10278 19369
rect 10220 19329 10232 19363
rect 10266 19360 10278 19363
rect 10594 19360 10600 19372
rect 10266 19332 10600 19360
rect 10266 19329 10278 19332
rect 10220 19323 10278 19329
rect 10594 19320 10600 19332
rect 10652 19320 10658 19372
rect 11514 19320 11520 19372
rect 11572 19320 11578 19372
rect 11716 19360 11744 19468
rect 12066 19456 12072 19508
rect 12124 19456 12130 19508
rect 12894 19496 12900 19508
rect 12452 19468 12900 19496
rect 11784 19431 11842 19437
rect 11784 19397 11796 19431
rect 11830 19428 11842 19431
rect 12084 19428 12112 19456
rect 12452 19440 12480 19468
rect 12894 19456 12900 19468
rect 12952 19456 12958 19508
rect 18601 19499 18659 19505
rect 18601 19465 18613 19499
rect 18647 19496 18659 19499
rect 18966 19496 18972 19508
rect 18647 19468 18972 19496
rect 18647 19465 18659 19468
rect 18601 19459 18659 19465
rect 18966 19456 18972 19468
rect 19024 19456 19030 19508
rect 19245 19499 19303 19505
rect 19245 19465 19257 19499
rect 19291 19465 19303 19499
rect 19245 19459 19303 19465
rect 19613 19499 19671 19505
rect 19613 19465 19625 19499
rect 19659 19496 19671 19499
rect 20162 19496 20168 19508
rect 19659 19468 20168 19496
rect 19659 19465 19671 19468
rect 19613 19459 19671 19465
rect 11830 19400 12112 19428
rect 11830 19397 11842 19400
rect 11784 19391 11842 19397
rect 12434 19388 12440 19440
rect 12492 19388 12498 19440
rect 14366 19388 14372 19440
rect 14424 19428 14430 19440
rect 14642 19428 14648 19440
rect 14424 19400 14648 19428
rect 14424 19388 14430 19400
rect 14642 19388 14648 19400
rect 14700 19428 14706 19440
rect 14921 19431 14979 19437
rect 14700 19400 14872 19428
rect 14700 19388 14706 19400
rect 12158 19360 12164 19372
rect 11716 19332 12164 19360
rect 12158 19320 12164 19332
rect 12216 19320 12222 19372
rect 14844 19369 14872 19400
rect 14921 19397 14933 19431
rect 14967 19428 14979 19431
rect 15930 19428 15936 19440
rect 14967 19400 15936 19428
rect 14967 19397 14979 19400
rect 14921 19391 14979 19397
rect 15930 19388 15936 19400
rect 15988 19388 15994 19440
rect 17494 19437 17500 19440
rect 17488 19428 17500 19437
rect 17455 19400 17500 19428
rect 17488 19391 17500 19400
rect 17494 19388 17500 19391
rect 17552 19388 17558 19440
rect 13357 19363 13415 19369
rect 13357 19329 13369 19363
rect 13403 19360 13415 19363
rect 13817 19363 13875 19369
rect 13817 19360 13829 19363
rect 13403 19332 13829 19360
rect 13403 19329 13415 19332
rect 13357 19323 13415 19329
rect 13817 19329 13829 19332
rect 13863 19329 13875 19363
rect 13817 19323 13875 19329
rect 14829 19363 14887 19369
rect 14829 19329 14841 19363
rect 14875 19329 14887 19363
rect 14829 19323 14887 19329
rect 15105 19363 15163 19369
rect 15105 19329 15117 19363
rect 15151 19329 15163 19363
rect 15105 19323 15163 19329
rect 17221 19363 17279 19369
rect 17221 19329 17233 19363
rect 17267 19360 17279 19363
rect 17310 19360 17316 19372
rect 17267 19332 17316 19360
rect 17267 19329 17279 19332
rect 17221 19323 17279 19329
rect 6196 19264 6500 19292
rect 6196 19233 6224 19264
rect 8202 19252 8208 19304
rect 8260 19252 8266 19304
rect 8294 19252 8300 19304
rect 8352 19252 8358 19304
rect 8389 19295 8447 19301
rect 8389 19261 8401 19295
rect 8435 19261 8447 19295
rect 8389 19255 8447 19261
rect 6181 19227 6239 19233
rect 6181 19193 6193 19227
rect 6227 19193 6239 19227
rect 6181 19187 6239 19193
rect 7742 19184 7748 19236
rect 7800 19184 7806 19236
rect 8220 19224 8248 19252
rect 8404 19224 8432 19255
rect 13446 19252 13452 19304
rect 13504 19252 13510 19304
rect 13633 19295 13691 19301
rect 13633 19261 13645 19295
rect 13679 19292 13691 19295
rect 13722 19292 13728 19304
rect 13679 19264 13728 19292
rect 13679 19261 13691 19264
rect 13633 19255 13691 19261
rect 13722 19252 13728 19264
rect 13780 19252 13786 19304
rect 14366 19252 14372 19304
rect 14424 19252 14430 19304
rect 15120 19224 15148 19323
rect 17310 19320 17316 19332
rect 17368 19360 17374 19372
rect 18877 19363 18935 19369
rect 17368 19332 18276 19360
rect 17368 19320 17374 19332
rect 18248 19292 18276 19332
rect 18877 19329 18889 19363
rect 18923 19360 18935 19363
rect 19260 19360 19288 19459
rect 20162 19456 20168 19468
rect 20220 19456 20226 19508
rect 20990 19456 20996 19508
rect 21048 19456 21054 19508
rect 21637 19499 21695 19505
rect 21637 19465 21649 19499
rect 21683 19496 21695 19499
rect 22094 19496 22100 19508
rect 21683 19468 22100 19496
rect 21683 19465 21695 19468
rect 21637 19459 21695 19465
rect 22094 19456 22100 19468
rect 22152 19456 22158 19508
rect 24854 19456 24860 19508
rect 24912 19496 24918 19508
rect 26973 19499 27031 19505
rect 26973 19496 26985 19499
rect 24912 19468 26985 19496
rect 24912 19456 24918 19468
rect 26973 19465 26985 19468
rect 27019 19465 27031 19499
rect 26973 19459 27031 19465
rect 20524 19431 20582 19437
rect 20524 19397 20536 19431
rect 20570 19428 20582 19431
rect 21008 19428 21036 19456
rect 27249 19431 27307 19437
rect 20570 19400 21036 19428
rect 23216 19400 26188 19428
rect 20570 19397 20582 19400
rect 20524 19391 20582 19397
rect 18923 19332 19288 19360
rect 18923 19329 18935 19332
rect 18877 19323 18935 19329
rect 19334 19320 19340 19372
rect 19392 19360 19398 19372
rect 19978 19360 19984 19372
rect 19392 19332 19984 19360
rect 19392 19320 19398 19332
rect 19978 19320 19984 19332
rect 20036 19360 20042 19372
rect 20257 19363 20315 19369
rect 20257 19360 20269 19363
rect 20036 19332 20269 19360
rect 20036 19320 20042 19332
rect 20257 19329 20269 19332
rect 20303 19329 20315 19363
rect 20257 19323 20315 19329
rect 22646 19320 22652 19372
rect 22704 19360 22710 19372
rect 23216 19369 23244 19400
rect 26160 19372 26188 19400
rect 27249 19397 27261 19431
rect 27295 19428 27307 19431
rect 27982 19428 27988 19440
rect 27295 19400 27988 19428
rect 27295 19397 27307 19400
rect 27249 19391 27307 19397
rect 27982 19388 27988 19400
rect 28040 19388 28046 19440
rect 22934 19363 22992 19369
rect 22934 19360 22946 19363
rect 22704 19332 22946 19360
rect 22704 19320 22710 19332
rect 22934 19329 22946 19332
rect 22980 19329 22992 19363
rect 22934 19323 22992 19329
rect 23201 19363 23259 19369
rect 23201 19329 23213 19363
rect 23247 19329 23259 19363
rect 23201 19323 23259 19329
rect 25958 19320 25964 19372
rect 26016 19320 26022 19372
rect 26142 19320 26148 19372
rect 26200 19320 26206 19372
rect 26418 19320 26424 19372
rect 26476 19320 26482 19372
rect 27152 19363 27210 19369
rect 27152 19329 27164 19363
rect 27198 19360 27210 19363
rect 27198 19332 27292 19360
rect 27198 19329 27210 19332
rect 27152 19323 27210 19329
rect 19352 19292 19380 19320
rect 18248 19264 19380 19292
rect 19702 19252 19708 19304
rect 19760 19252 19766 19304
rect 19889 19295 19947 19301
rect 19889 19261 19901 19295
rect 19935 19292 19947 19295
rect 20070 19292 20076 19304
rect 19935 19264 20076 19292
rect 19935 19261 19947 19264
rect 19889 19255 19947 19261
rect 20070 19252 20076 19264
rect 20128 19252 20134 19304
rect 27264 19292 27292 19332
rect 27338 19320 27344 19372
rect 27396 19320 27402 19372
rect 27522 19360 27528 19372
rect 27483 19332 27528 19360
rect 27522 19320 27528 19332
rect 27580 19320 27586 19372
rect 27617 19363 27675 19369
rect 27617 19329 27629 19363
rect 27663 19360 27675 19363
rect 29362 19360 29368 19372
rect 27663 19332 29368 19360
rect 27663 19329 27675 19332
rect 27617 19323 27675 19329
rect 29362 19320 29368 19332
rect 29420 19320 29426 19372
rect 28718 19292 28724 19304
rect 27264 19264 28724 19292
rect 28718 19252 28724 19264
rect 28776 19252 28782 19304
rect 8220 19196 8432 19224
rect 12820 19196 15148 19224
rect 5902 19116 5908 19168
rect 5960 19156 5966 19168
rect 12820 19156 12848 19196
rect 5960 19128 12848 19156
rect 5960 19116 5966 19128
rect 12986 19116 12992 19168
rect 13044 19116 13050 19168
rect 15286 19116 15292 19168
rect 15344 19116 15350 19168
rect 19061 19159 19119 19165
rect 19061 19125 19073 19159
rect 19107 19156 19119 19159
rect 19334 19156 19340 19168
rect 19107 19128 19340 19156
rect 19107 19125 19119 19128
rect 19061 19119 19119 19125
rect 19334 19116 19340 19128
rect 19392 19116 19398 19168
rect 21821 19159 21879 19165
rect 21821 19125 21833 19159
rect 21867 19156 21879 19159
rect 22830 19156 22836 19168
rect 21867 19128 22836 19156
rect 21867 19125 21879 19128
rect 21821 19119 21879 19125
rect 22830 19116 22836 19128
rect 22888 19116 22894 19168
rect 23014 19116 23020 19168
rect 23072 19156 23078 19168
rect 25222 19156 25228 19168
rect 23072 19128 25228 19156
rect 23072 19116 23078 19128
rect 25222 19116 25228 19128
rect 25280 19116 25286 19168
rect 25774 19116 25780 19168
rect 25832 19116 25838 19168
rect 26602 19116 26608 19168
rect 26660 19116 26666 19168
rect 29454 19116 29460 19168
rect 29512 19156 29518 19168
rect 30650 19156 30656 19168
rect 29512 19128 30656 19156
rect 29512 19116 29518 19128
rect 30650 19116 30656 19128
rect 30708 19116 30714 19168
rect 1104 19066 31832 19088
rect 1104 19014 4182 19066
rect 4234 19014 4246 19066
rect 4298 19014 4310 19066
rect 4362 19014 4374 19066
rect 4426 19014 4438 19066
rect 4490 19014 4502 19066
rect 4554 19014 10182 19066
rect 10234 19014 10246 19066
rect 10298 19014 10310 19066
rect 10362 19014 10374 19066
rect 10426 19014 10438 19066
rect 10490 19014 10502 19066
rect 10554 19014 16182 19066
rect 16234 19014 16246 19066
rect 16298 19014 16310 19066
rect 16362 19014 16374 19066
rect 16426 19014 16438 19066
rect 16490 19014 16502 19066
rect 16554 19014 22182 19066
rect 22234 19014 22246 19066
rect 22298 19014 22310 19066
rect 22362 19014 22374 19066
rect 22426 19014 22438 19066
rect 22490 19014 22502 19066
rect 22554 19014 28182 19066
rect 28234 19014 28246 19066
rect 28298 19014 28310 19066
rect 28362 19014 28374 19066
rect 28426 19014 28438 19066
rect 28490 19014 28502 19066
rect 28554 19014 31832 19066
rect 1104 18992 31832 19014
rect 3050 18912 3056 18964
rect 3108 18912 3114 18964
rect 4062 18912 4068 18964
rect 4120 18912 4126 18964
rect 5534 18912 5540 18964
rect 5592 18912 5598 18964
rect 5902 18912 5908 18964
rect 5960 18912 5966 18964
rect 5994 18912 6000 18964
rect 6052 18952 6058 18964
rect 6641 18955 6699 18961
rect 6641 18952 6653 18955
rect 6052 18924 6653 18952
rect 6052 18912 6058 18924
rect 6641 18921 6653 18924
rect 6687 18921 6699 18955
rect 6641 18915 6699 18921
rect 10594 18912 10600 18964
rect 10652 18912 10658 18964
rect 11606 18952 11612 18964
rect 10796 18924 11612 18952
rect 2961 18887 3019 18893
rect 2961 18853 2973 18887
rect 3007 18884 3019 18887
rect 4080 18884 4108 18912
rect 3007 18856 4108 18884
rect 3007 18853 3019 18856
rect 2961 18847 3019 18853
rect 4433 18819 4491 18825
rect 4433 18785 4445 18819
rect 4479 18816 4491 18819
rect 4614 18816 4620 18828
rect 4479 18788 4620 18816
rect 4479 18785 4491 18788
rect 4433 18779 4491 18785
rect 4614 18776 4620 18788
rect 4672 18776 4678 18828
rect 5166 18776 5172 18828
rect 5224 18776 5230 18828
rect 934 18708 940 18760
rect 992 18748 998 18760
rect 1397 18751 1455 18757
rect 1397 18748 1409 18751
rect 992 18720 1409 18748
rect 992 18708 998 18720
rect 1397 18717 1409 18720
rect 1443 18717 1455 18751
rect 1397 18711 1455 18717
rect 2777 18751 2835 18757
rect 2777 18717 2789 18751
rect 2823 18748 2835 18751
rect 3142 18748 3148 18760
rect 2823 18720 3148 18748
rect 2823 18717 2835 18720
rect 2777 18711 2835 18717
rect 3142 18708 3148 18720
rect 3200 18708 3206 18760
rect 3237 18751 3295 18757
rect 3237 18717 3249 18751
rect 3283 18748 3295 18751
rect 5184 18748 5212 18776
rect 5353 18751 5411 18757
rect 5353 18748 5365 18751
rect 3283 18720 3832 18748
rect 5184 18720 5365 18748
rect 3283 18717 3295 18720
rect 3237 18711 3295 18717
rect 1581 18615 1639 18621
rect 1581 18581 1593 18615
rect 1627 18612 1639 18615
rect 3694 18612 3700 18624
rect 1627 18584 3700 18612
rect 1627 18581 1639 18584
rect 1581 18575 1639 18581
rect 3694 18572 3700 18584
rect 3752 18572 3758 18624
rect 3804 18621 3832 18720
rect 5353 18717 5365 18720
rect 5399 18717 5411 18751
rect 5552 18748 5580 18912
rect 10796 18884 10824 18924
rect 7300 18856 10824 18884
rect 10873 18887 10931 18893
rect 7098 18776 7104 18828
rect 7156 18776 7162 18828
rect 7190 18776 7196 18828
rect 7248 18816 7254 18828
rect 7300 18825 7328 18856
rect 10873 18853 10885 18887
rect 10919 18853 10931 18887
rect 10873 18847 10931 18853
rect 7285 18819 7343 18825
rect 7285 18816 7297 18819
rect 7248 18788 7297 18816
rect 7248 18776 7254 18788
rect 7285 18785 7297 18788
rect 7331 18785 7343 18819
rect 7285 18779 7343 18785
rect 7742 18776 7748 18828
rect 7800 18816 7806 18828
rect 8021 18819 8079 18825
rect 8021 18816 8033 18819
rect 7800 18788 8033 18816
rect 7800 18776 7806 18788
rect 8021 18785 8033 18788
rect 8067 18785 8079 18819
rect 8021 18779 8079 18785
rect 5629 18751 5687 18757
rect 5629 18748 5641 18751
rect 5552 18720 5641 18748
rect 5353 18711 5411 18717
rect 5629 18717 5641 18720
rect 5675 18717 5687 18751
rect 5629 18711 5687 18717
rect 5721 18751 5779 18757
rect 5721 18717 5733 18751
rect 5767 18748 5779 18751
rect 5810 18748 5816 18760
rect 5767 18720 5816 18748
rect 5767 18717 5779 18720
rect 5721 18711 5779 18717
rect 5810 18708 5816 18720
rect 5868 18708 5874 18760
rect 10781 18751 10839 18757
rect 10781 18717 10793 18751
rect 10827 18748 10839 18751
rect 10888 18748 10916 18847
rect 11440 18825 11468 18924
rect 11606 18912 11612 18924
rect 11664 18952 11670 18964
rect 11974 18952 11980 18964
rect 11664 18924 11980 18952
rect 11664 18912 11670 18924
rect 11974 18912 11980 18924
rect 12032 18912 12038 18964
rect 13173 18955 13231 18961
rect 13173 18921 13185 18955
rect 13219 18952 13231 18955
rect 14366 18952 14372 18964
rect 13219 18924 14372 18952
rect 13219 18921 13231 18924
rect 13173 18915 13231 18921
rect 11425 18819 11483 18825
rect 11425 18785 11437 18819
rect 11471 18785 11483 18819
rect 11425 18779 11483 18785
rect 11514 18776 11520 18828
rect 11572 18816 11578 18828
rect 11793 18819 11851 18825
rect 11793 18816 11805 18819
rect 11572 18788 11805 18816
rect 11572 18776 11578 18788
rect 11793 18785 11805 18788
rect 11839 18785 11851 18819
rect 11793 18779 11851 18785
rect 10827 18720 10916 18748
rect 11241 18751 11299 18757
rect 10827 18717 10839 18720
rect 10781 18711 10839 18717
rect 11241 18717 11253 18751
rect 11287 18748 11299 18751
rect 11330 18748 11336 18760
rect 11287 18720 11336 18748
rect 11287 18717 11299 18720
rect 11241 18711 11299 18717
rect 11330 18708 11336 18720
rect 11388 18708 11394 18760
rect 13262 18708 13268 18760
rect 13320 18708 13326 18760
rect 13372 18757 13400 18924
rect 14366 18912 14372 18924
rect 14424 18912 14430 18964
rect 15378 18952 15384 18964
rect 14752 18924 15384 18952
rect 13909 18887 13967 18893
rect 13909 18853 13921 18887
rect 13955 18884 13967 18887
rect 14752 18884 14780 18924
rect 15378 18912 15384 18924
rect 15436 18912 15442 18964
rect 15930 18912 15936 18964
rect 15988 18952 15994 18964
rect 16117 18955 16175 18961
rect 16117 18952 16129 18955
rect 15988 18924 16129 18952
rect 15988 18912 15994 18924
rect 16117 18921 16129 18924
rect 16163 18921 16175 18955
rect 16117 18915 16175 18921
rect 17589 18955 17647 18961
rect 17589 18921 17601 18955
rect 17635 18952 17647 18955
rect 17678 18952 17684 18964
rect 17635 18924 17684 18952
rect 17635 18921 17647 18924
rect 17589 18915 17647 18921
rect 13955 18856 14780 18884
rect 13955 18853 13967 18856
rect 13909 18847 13967 18853
rect 16132 18816 16160 18915
rect 17678 18912 17684 18924
rect 17736 18912 17742 18964
rect 19610 18952 19616 18964
rect 17880 18924 19616 18952
rect 16666 18844 16672 18896
rect 16724 18884 16730 18896
rect 17129 18887 17187 18893
rect 17129 18884 17141 18887
rect 16724 18856 17141 18884
rect 16724 18844 16730 18856
rect 17129 18853 17141 18856
rect 17175 18853 17187 18887
rect 17129 18847 17187 18853
rect 16761 18819 16819 18825
rect 16761 18816 16773 18819
rect 13464 18788 14872 18816
rect 16132 18788 16773 18816
rect 13358 18751 13416 18757
rect 13358 18717 13370 18751
rect 13404 18717 13416 18751
rect 13358 18711 13416 18717
rect 4157 18683 4215 18689
rect 4157 18649 4169 18683
rect 4203 18680 4215 18683
rect 4617 18683 4675 18689
rect 4617 18680 4629 18683
rect 4203 18652 4629 18680
rect 4203 18649 4215 18652
rect 4157 18643 4215 18649
rect 4617 18649 4629 18652
rect 4663 18649 4675 18683
rect 4617 18643 4675 18649
rect 5534 18640 5540 18692
rect 5592 18640 5598 18692
rect 7009 18683 7067 18689
rect 7009 18649 7021 18683
rect 7055 18680 7067 18683
rect 7469 18683 7527 18689
rect 7469 18680 7481 18683
rect 7055 18652 7481 18680
rect 7055 18649 7067 18652
rect 7009 18643 7067 18649
rect 7469 18649 7481 18652
rect 7515 18649 7527 18683
rect 7469 18643 7527 18649
rect 11882 18640 11888 18692
rect 11940 18680 11946 18692
rect 12038 18683 12096 18689
rect 12038 18680 12050 18683
rect 11940 18652 12050 18680
rect 11940 18640 11946 18652
rect 12038 18649 12050 18652
rect 12084 18649 12096 18683
rect 12038 18643 12096 18649
rect 13464 18624 13492 18788
rect 13771 18751 13829 18757
rect 13771 18717 13783 18751
rect 13817 18748 13829 18751
rect 14182 18748 14188 18760
rect 13817 18720 14188 18748
rect 13817 18717 13829 18720
rect 13771 18711 13829 18717
rect 14182 18708 14188 18720
rect 14240 18708 14246 18760
rect 14274 18708 14280 18760
rect 14332 18708 14338 18760
rect 14458 18708 14464 18760
rect 14516 18708 14522 18760
rect 14550 18708 14556 18760
rect 14608 18748 14614 18760
rect 14737 18751 14795 18757
rect 14737 18748 14749 18751
rect 14608 18720 14749 18748
rect 14608 18708 14614 18720
rect 14737 18717 14749 18720
rect 14783 18717 14795 18751
rect 14844 18748 14872 18788
rect 16761 18785 16773 18788
rect 16807 18785 16819 18819
rect 17144 18816 17172 18847
rect 17880 18816 17908 18924
rect 19610 18912 19616 18924
rect 19668 18912 19674 18964
rect 20625 18955 20683 18961
rect 20625 18921 20637 18955
rect 20671 18952 20683 18955
rect 20714 18952 20720 18964
rect 20671 18924 20720 18952
rect 20671 18921 20683 18924
rect 20625 18915 20683 18921
rect 20714 18912 20720 18924
rect 20772 18912 20778 18964
rect 21174 18912 21180 18964
rect 21232 18912 21238 18964
rect 27982 18912 27988 18964
rect 28040 18952 28046 18964
rect 28353 18955 28411 18961
rect 28353 18952 28365 18955
rect 28040 18924 28365 18952
rect 28040 18912 28046 18924
rect 28353 18921 28365 18924
rect 28399 18921 28411 18955
rect 28353 18915 28411 18921
rect 19242 18844 19248 18896
rect 19300 18844 19306 18896
rect 21085 18887 21143 18893
rect 21085 18853 21097 18887
rect 21131 18884 21143 18887
rect 22462 18884 22468 18896
rect 21131 18856 22468 18884
rect 21131 18853 21143 18856
rect 21085 18847 21143 18853
rect 22462 18844 22468 18856
rect 22520 18844 22526 18896
rect 22572 18856 23152 18884
rect 17144 18788 17908 18816
rect 16761 18779 16819 18785
rect 18230 18776 18236 18828
rect 18288 18776 18294 18828
rect 16945 18751 17003 18757
rect 16945 18748 16957 18751
rect 14844 18720 16957 18748
rect 14737 18711 14795 18717
rect 16945 18717 16957 18720
rect 16991 18717 17003 18751
rect 16945 18711 17003 18717
rect 17957 18751 18015 18757
rect 17957 18717 17969 18751
rect 18003 18748 18015 18751
rect 18322 18748 18328 18760
rect 18003 18720 18328 18748
rect 18003 18717 18015 18720
rect 17957 18711 18015 18717
rect 13541 18683 13599 18689
rect 13541 18649 13553 18683
rect 13587 18649 13599 18683
rect 13541 18643 13599 18649
rect 13633 18683 13691 18689
rect 13633 18649 13645 18683
rect 13679 18680 13691 18683
rect 13906 18680 13912 18692
rect 13679 18652 13912 18680
rect 13679 18649 13691 18652
rect 13633 18643 13691 18649
rect 3789 18615 3847 18621
rect 3789 18581 3801 18615
rect 3835 18581 3847 18615
rect 3789 18575 3847 18581
rect 4249 18615 4307 18621
rect 4249 18581 4261 18615
rect 4295 18612 4307 18615
rect 4798 18612 4804 18624
rect 4295 18584 4804 18612
rect 4295 18581 4307 18584
rect 4249 18575 4307 18581
rect 4798 18572 4804 18584
rect 4856 18612 4862 18624
rect 7558 18612 7564 18624
rect 4856 18584 7564 18612
rect 4856 18572 4862 18584
rect 7558 18572 7564 18584
rect 7616 18612 7622 18624
rect 11333 18615 11391 18621
rect 11333 18612 11345 18615
rect 7616 18584 11345 18612
rect 7616 18572 7622 18584
rect 11333 18581 11345 18584
rect 11379 18612 11391 18615
rect 13446 18612 13452 18624
rect 11379 18584 13452 18612
rect 11379 18581 11391 18584
rect 11333 18575 11391 18581
rect 13446 18572 13452 18584
rect 13504 18572 13510 18624
rect 13556 18612 13584 18643
rect 13906 18640 13912 18652
rect 13964 18640 13970 18692
rect 13814 18612 13820 18624
rect 13556 18584 13820 18612
rect 13814 18572 13820 18584
rect 13872 18612 13878 18624
rect 14292 18612 14320 18708
rect 14982 18683 15040 18689
rect 14982 18680 14994 18683
rect 14660 18652 14994 18680
rect 14660 18621 14688 18652
rect 14982 18649 14994 18652
rect 15028 18649 15040 18683
rect 16960 18680 16988 18711
rect 18322 18708 18328 18720
rect 18380 18708 18386 18760
rect 19260 18757 19288 18844
rect 21634 18776 21640 18828
rect 21692 18776 21698 18828
rect 21821 18819 21879 18825
rect 21821 18785 21833 18819
rect 21867 18785 21879 18819
rect 21821 18779 21879 18785
rect 18509 18751 18567 18757
rect 18509 18717 18521 18751
rect 18555 18748 18567 18751
rect 19245 18751 19303 18757
rect 18555 18720 19196 18748
rect 18555 18717 18567 18720
rect 18509 18711 18567 18717
rect 18046 18680 18052 18692
rect 16960 18652 18052 18680
rect 14982 18643 15040 18649
rect 18046 18640 18052 18652
rect 18104 18640 18110 18692
rect 13872 18584 14320 18612
rect 14645 18615 14703 18621
rect 13872 18572 13878 18584
rect 14645 18581 14657 18615
rect 14691 18581 14703 18615
rect 14645 18575 14703 18581
rect 16206 18572 16212 18624
rect 16264 18572 16270 18624
rect 19058 18572 19064 18624
rect 19116 18572 19122 18624
rect 19168 18612 19196 18720
rect 19245 18717 19257 18751
rect 19291 18717 19303 18751
rect 19245 18711 19303 18717
rect 20901 18751 20959 18757
rect 20901 18717 20913 18751
rect 20947 18748 20959 18751
rect 21450 18748 21456 18760
rect 20947 18720 21456 18748
rect 20947 18717 20959 18720
rect 20901 18711 20959 18717
rect 21450 18708 21456 18720
rect 21508 18708 21514 18760
rect 21836 18748 21864 18779
rect 22094 18776 22100 18828
rect 22152 18816 22158 18828
rect 22572 18825 22600 18856
rect 22557 18819 22615 18825
rect 22557 18816 22569 18819
rect 22152 18788 22569 18816
rect 22152 18776 22158 18788
rect 22557 18785 22569 18788
rect 22603 18785 22615 18819
rect 23014 18816 23020 18828
rect 22557 18779 22615 18785
rect 22664 18788 23020 18816
rect 22664 18748 22692 18788
rect 23014 18776 23020 18788
rect 23072 18776 23078 18828
rect 23124 18816 23152 18856
rect 23124 18788 23336 18816
rect 21836 18720 22692 18748
rect 22925 18751 22983 18757
rect 22925 18717 22937 18751
rect 22971 18748 22983 18751
rect 23198 18748 23204 18760
rect 22971 18720 23204 18748
rect 22971 18717 22983 18720
rect 22925 18711 22983 18717
rect 19334 18640 19340 18692
rect 19392 18680 19398 18692
rect 19490 18683 19548 18689
rect 19490 18680 19502 18683
rect 19392 18652 19502 18680
rect 19392 18640 19398 18652
rect 19490 18649 19502 18652
rect 19536 18649 19548 18683
rect 19490 18643 19548 18649
rect 21545 18683 21603 18689
rect 21545 18649 21557 18683
rect 21591 18680 21603 18683
rect 22005 18683 22063 18689
rect 22005 18680 22017 18683
rect 21591 18652 22017 18680
rect 21591 18649 21603 18652
rect 21545 18643 21603 18649
rect 22005 18649 22017 18652
rect 22051 18649 22063 18683
rect 22005 18643 22063 18649
rect 19610 18612 19616 18624
rect 19168 18584 19616 18612
rect 19610 18572 19616 18584
rect 19668 18572 19674 18624
rect 22738 18572 22744 18624
rect 22796 18572 22802 18624
rect 22830 18572 22836 18624
rect 22888 18612 22894 18624
rect 22940 18612 22968 18711
rect 23198 18708 23204 18720
rect 23256 18708 23262 18760
rect 23308 18757 23336 18788
rect 23293 18751 23351 18757
rect 23293 18717 23305 18751
rect 23339 18717 23351 18751
rect 23293 18711 23351 18717
rect 25501 18751 25559 18757
rect 25501 18717 25513 18751
rect 25547 18748 25559 18751
rect 26142 18748 26148 18760
rect 25547 18720 26148 18748
rect 25547 18717 25559 18720
rect 25501 18711 25559 18717
rect 26142 18708 26148 18720
rect 26200 18748 26206 18760
rect 26973 18751 27031 18757
rect 26973 18748 26985 18751
rect 26200 18720 26985 18748
rect 26200 18708 26206 18720
rect 26973 18717 26985 18720
rect 27019 18748 27031 18751
rect 27019 18720 27384 18748
rect 27019 18717 27031 18720
rect 26973 18711 27031 18717
rect 23014 18640 23020 18692
rect 23072 18640 23078 18692
rect 23109 18683 23167 18689
rect 23109 18649 23121 18683
rect 23155 18680 23167 18683
rect 23382 18680 23388 18692
rect 23155 18652 23388 18680
rect 23155 18649 23167 18652
rect 23109 18643 23167 18649
rect 23382 18640 23388 18652
rect 23440 18640 23446 18692
rect 25774 18689 25780 18692
rect 25768 18680 25780 18689
rect 25735 18652 25780 18680
rect 25768 18643 25780 18652
rect 25774 18640 25780 18643
rect 25832 18640 25838 18692
rect 26602 18640 26608 18692
rect 26660 18680 26666 18692
rect 27218 18683 27276 18689
rect 27218 18680 27230 18683
rect 26660 18652 27230 18680
rect 26660 18640 26666 18652
rect 27218 18649 27230 18652
rect 27264 18649 27276 18683
rect 27356 18680 27384 18720
rect 27522 18708 27528 18760
rect 27580 18748 27586 18760
rect 28997 18751 29055 18757
rect 28997 18748 29009 18751
rect 27580 18720 29009 18748
rect 27580 18708 27586 18720
rect 28997 18717 29009 18720
rect 29043 18717 29055 18751
rect 28997 18711 29055 18717
rect 30558 18680 30564 18692
rect 27356 18652 30564 18680
rect 27218 18643 27276 18649
rect 30558 18640 30564 18652
rect 30616 18640 30622 18692
rect 22888 18584 22968 18612
rect 26881 18615 26939 18621
rect 22888 18572 22894 18584
rect 26881 18581 26893 18615
rect 26927 18612 26939 18615
rect 27522 18612 27528 18624
rect 26927 18584 27528 18612
rect 26927 18581 26939 18584
rect 26881 18575 26939 18581
rect 27522 18572 27528 18584
rect 27580 18572 27586 18624
rect 28442 18572 28448 18624
rect 28500 18572 28506 18624
rect 1104 18522 31832 18544
rect 1104 18470 4922 18522
rect 4974 18470 4986 18522
rect 5038 18470 5050 18522
rect 5102 18470 5114 18522
rect 5166 18470 5178 18522
rect 5230 18470 5242 18522
rect 5294 18470 10922 18522
rect 10974 18470 10986 18522
rect 11038 18470 11050 18522
rect 11102 18470 11114 18522
rect 11166 18470 11178 18522
rect 11230 18470 11242 18522
rect 11294 18470 16922 18522
rect 16974 18470 16986 18522
rect 17038 18470 17050 18522
rect 17102 18470 17114 18522
rect 17166 18470 17178 18522
rect 17230 18470 17242 18522
rect 17294 18470 22922 18522
rect 22974 18470 22986 18522
rect 23038 18470 23050 18522
rect 23102 18470 23114 18522
rect 23166 18470 23178 18522
rect 23230 18470 23242 18522
rect 23294 18470 28922 18522
rect 28974 18470 28986 18522
rect 29038 18470 29050 18522
rect 29102 18470 29114 18522
rect 29166 18470 29178 18522
rect 29230 18470 29242 18522
rect 29294 18470 31832 18522
rect 1104 18448 31832 18470
rect 7837 18411 7895 18417
rect 7837 18377 7849 18411
rect 7883 18377 7895 18411
rect 7837 18371 7895 18377
rect 7653 18275 7711 18281
rect 7653 18241 7665 18275
rect 7699 18272 7711 18275
rect 7852 18272 7880 18371
rect 11882 18368 11888 18420
rect 11940 18368 11946 18420
rect 12161 18411 12219 18417
rect 12161 18377 12173 18411
rect 12207 18408 12219 18411
rect 12250 18408 12256 18420
rect 12207 18380 12256 18408
rect 12207 18377 12219 18380
rect 12161 18371 12219 18377
rect 12250 18368 12256 18380
rect 12308 18368 12314 18420
rect 12529 18411 12587 18417
rect 12529 18377 12541 18411
rect 12575 18408 12587 18411
rect 12802 18408 12808 18420
rect 12575 18380 12808 18408
rect 12575 18377 12587 18380
rect 12529 18371 12587 18377
rect 12802 18368 12808 18380
rect 12860 18368 12866 18420
rect 12894 18368 12900 18420
rect 12952 18408 12958 18420
rect 13170 18408 13176 18420
rect 12952 18380 13176 18408
rect 12952 18368 12958 18380
rect 13170 18368 13176 18380
rect 13228 18408 13234 18420
rect 14090 18408 14096 18420
rect 13228 18380 14096 18408
rect 13228 18368 13234 18380
rect 14090 18368 14096 18380
rect 14148 18368 14154 18420
rect 14458 18368 14464 18420
rect 14516 18408 14522 18420
rect 15105 18411 15163 18417
rect 15105 18408 15117 18411
rect 14516 18380 15117 18408
rect 14516 18368 14522 18380
rect 15105 18377 15117 18380
rect 15151 18377 15163 18411
rect 15105 18371 15163 18377
rect 15473 18411 15531 18417
rect 15473 18377 15485 18411
rect 15519 18408 15531 18411
rect 16206 18408 16212 18420
rect 15519 18380 16212 18408
rect 15519 18377 15531 18380
rect 15473 18371 15531 18377
rect 16206 18368 16212 18380
rect 16264 18368 16270 18420
rect 16666 18368 16672 18420
rect 16724 18368 16730 18420
rect 17221 18411 17279 18417
rect 17221 18377 17233 18411
rect 17267 18377 17279 18411
rect 17221 18371 17279 18377
rect 12621 18343 12679 18349
rect 12621 18309 12633 18343
rect 12667 18340 12679 18343
rect 15010 18340 15016 18352
rect 12667 18312 15016 18340
rect 12667 18309 12679 18312
rect 12621 18303 12679 18309
rect 15010 18300 15016 18312
rect 15068 18340 15074 18352
rect 15565 18343 15623 18349
rect 15565 18340 15577 18343
rect 15068 18312 15577 18340
rect 15068 18300 15074 18312
rect 15565 18309 15577 18312
rect 15611 18340 15623 18343
rect 16684 18340 16712 18368
rect 15611 18312 16712 18340
rect 17236 18340 17264 18371
rect 18046 18368 18052 18420
rect 18104 18368 18110 18420
rect 19058 18368 19064 18420
rect 19116 18408 19122 18420
rect 19153 18411 19211 18417
rect 19153 18408 19165 18411
rect 19116 18380 19165 18408
rect 19116 18368 19122 18380
rect 19153 18377 19165 18380
rect 19199 18377 19211 18411
rect 19153 18371 19211 18377
rect 19334 18368 19340 18420
rect 19392 18408 19398 18420
rect 21637 18411 21695 18417
rect 21637 18408 21649 18411
rect 19392 18380 21649 18408
rect 19392 18368 19398 18380
rect 21637 18377 21649 18380
rect 21683 18377 21695 18411
rect 21637 18371 21695 18377
rect 21726 18368 21732 18420
rect 21784 18368 21790 18420
rect 25958 18368 25964 18420
rect 26016 18368 26022 18420
rect 26329 18411 26387 18417
rect 26329 18377 26341 18411
rect 26375 18408 26387 18411
rect 28442 18408 28448 18420
rect 26375 18380 28448 18408
rect 26375 18377 26387 18380
rect 26329 18371 26387 18377
rect 28442 18368 28448 18380
rect 28500 18368 28506 18420
rect 17558 18343 17616 18349
rect 17558 18340 17570 18343
rect 17236 18312 17570 18340
rect 15611 18309 15623 18312
rect 15565 18303 15623 18309
rect 17558 18309 17570 18312
rect 17604 18309 17616 18343
rect 18064 18340 18092 18368
rect 19245 18343 19303 18349
rect 19245 18340 19257 18343
rect 18064 18312 19257 18340
rect 17558 18303 17616 18309
rect 19245 18309 19257 18312
rect 19291 18309 19303 18343
rect 19245 18303 19303 18309
rect 19702 18300 19708 18352
rect 19760 18340 19766 18352
rect 20073 18343 20131 18349
rect 20073 18340 20085 18343
rect 19760 18312 20085 18340
rect 19760 18300 19766 18312
rect 20073 18309 20085 18312
rect 20119 18340 20131 18343
rect 21744 18340 21772 18368
rect 28074 18340 28080 18352
rect 20119 18312 21772 18340
rect 26620 18312 28080 18340
rect 20119 18309 20131 18312
rect 20073 18303 20131 18309
rect 7699 18244 7880 18272
rect 8205 18275 8263 18281
rect 7699 18241 7711 18244
rect 7653 18235 7711 18241
rect 8205 18241 8217 18275
rect 8251 18272 8263 18275
rect 8665 18275 8723 18281
rect 8665 18272 8677 18275
rect 8251 18244 8677 18272
rect 8251 18241 8263 18244
rect 8205 18235 8263 18241
rect 8665 18241 8677 18244
rect 8711 18241 8723 18275
rect 8665 18235 8723 18241
rect 12069 18275 12127 18281
rect 12069 18241 12081 18275
rect 12115 18272 12127 18275
rect 12986 18272 12992 18284
rect 12115 18244 12992 18272
rect 12115 18241 12127 18244
rect 12069 18235 12127 18241
rect 12986 18232 12992 18244
rect 13044 18232 13050 18284
rect 13814 18272 13820 18284
rect 13096 18244 13820 18272
rect 8110 18164 8116 18216
rect 8168 18204 8174 18216
rect 8297 18207 8355 18213
rect 8297 18204 8309 18207
rect 8168 18176 8309 18204
rect 8168 18164 8174 18176
rect 8297 18173 8309 18176
rect 8343 18173 8355 18207
rect 8297 18167 8355 18173
rect 8478 18164 8484 18216
rect 8536 18164 8542 18216
rect 9214 18164 9220 18216
rect 9272 18164 9278 18216
rect 12805 18207 12863 18213
rect 12805 18204 12817 18207
rect 12406 18176 12817 18204
rect 8202 18096 8208 18148
rect 8260 18136 8266 18148
rect 12406 18136 12434 18176
rect 12805 18173 12817 18176
rect 12851 18204 12863 18207
rect 12894 18204 12900 18216
rect 12851 18176 12900 18204
rect 12851 18173 12863 18176
rect 12805 18167 12863 18173
rect 12894 18164 12900 18176
rect 12952 18164 12958 18216
rect 8260 18108 12434 18136
rect 8260 18096 8266 18108
rect 7282 18028 7288 18080
rect 7340 18068 7346 18080
rect 7469 18071 7527 18077
rect 7469 18068 7481 18071
rect 7340 18040 7481 18068
rect 7340 18028 7346 18040
rect 7469 18037 7481 18040
rect 7515 18037 7527 18071
rect 7469 18031 7527 18037
rect 9490 18028 9496 18080
rect 9548 18068 9554 18080
rect 13096 18068 13124 18244
rect 13814 18232 13820 18244
rect 13872 18232 13878 18284
rect 14274 18232 14280 18284
rect 14332 18281 14338 18284
rect 14332 18235 14344 18281
rect 17037 18275 17095 18281
rect 17037 18241 17049 18275
rect 17083 18241 17095 18275
rect 17037 18235 17095 18241
rect 14332 18232 14338 18235
rect 14550 18164 14556 18216
rect 14608 18164 14614 18216
rect 15654 18164 15660 18216
rect 15712 18164 15718 18216
rect 17052 18204 17080 18235
rect 17310 18232 17316 18284
rect 17368 18232 17374 18284
rect 19981 18275 20039 18281
rect 17420 18244 18828 18272
rect 17420 18204 17448 18244
rect 17052 18176 17448 18204
rect 9548 18040 13124 18068
rect 13173 18071 13231 18077
rect 9548 18028 9554 18040
rect 13173 18037 13185 18071
rect 13219 18068 13231 18071
rect 13906 18068 13912 18080
rect 13219 18040 13912 18068
rect 13219 18037 13231 18040
rect 13173 18031 13231 18037
rect 13906 18028 13912 18040
rect 13964 18028 13970 18080
rect 14182 18028 14188 18080
rect 14240 18068 14246 18080
rect 14568 18068 14596 18164
rect 18800 18145 18828 18244
rect 19981 18241 19993 18275
rect 20027 18272 20039 18275
rect 20441 18275 20499 18281
rect 20441 18272 20453 18275
rect 20027 18244 20453 18272
rect 20027 18241 20039 18244
rect 19981 18235 20039 18241
rect 20441 18241 20453 18244
rect 20487 18241 20499 18275
rect 20441 18235 20499 18241
rect 21174 18232 21180 18284
rect 21232 18232 21238 18284
rect 21453 18275 21511 18281
rect 21453 18241 21465 18275
rect 21499 18272 21511 18275
rect 24854 18272 24860 18284
rect 21499 18244 24860 18272
rect 21499 18241 21511 18244
rect 21453 18235 21511 18241
rect 24854 18232 24860 18244
rect 24912 18232 24918 18284
rect 19150 18164 19156 18216
rect 19208 18204 19214 18216
rect 19337 18207 19395 18213
rect 19337 18204 19349 18207
rect 19208 18176 19349 18204
rect 19208 18164 19214 18176
rect 19337 18173 19349 18176
rect 19383 18173 19395 18207
rect 19337 18167 19395 18173
rect 20254 18164 20260 18216
rect 20312 18164 20318 18216
rect 20346 18164 20352 18216
rect 20404 18204 20410 18216
rect 20993 18207 21051 18213
rect 20993 18204 21005 18207
rect 20404 18176 21005 18204
rect 20404 18164 20410 18176
rect 20993 18173 21005 18176
rect 21039 18173 21051 18207
rect 20993 18167 21051 18173
rect 21266 18164 21272 18216
rect 21324 18164 21330 18216
rect 22738 18204 22744 18216
rect 21468 18176 22744 18204
rect 18785 18139 18843 18145
rect 18785 18105 18797 18139
rect 18831 18105 18843 18139
rect 19518 18136 19524 18148
rect 18785 18099 18843 18105
rect 18892 18108 19524 18136
rect 14240 18040 14596 18068
rect 18693 18071 18751 18077
rect 14240 18028 14246 18040
rect 18693 18037 18705 18071
rect 18739 18068 18751 18071
rect 18892 18068 18920 18108
rect 19518 18096 19524 18108
rect 19576 18096 19582 18148
rect 18739 18040 18920 18068
rect 18739 18037 18751 18040
rect 18693 18031 18751 18037
rect 18966 18028 18972 18080
rect 19024 18068 19030 18080
rect 19613 18071 19671 18077
rect 19613 18068 19625 18071
rect 19024 18040 19625 18068
rect 19024 18028 19030 18040
rect 19613 18037 19625 18040
rect 19659 18037 19671 18071
rect 19613 18031 19671 18037
rect 20070 18028 20076 18080
rect 20128 18068 20134 18080
rect 20806 18068 20812 18080
rect 20128 18040 20812 18068
rect 20128 18028 20134 18040
rect 20806 18028 20812 18040
rect 20864 18028 20870 18080
rect 21468 18077 21496 18176
rect 22738 18164 22744 18176
rect 22796 18164 22802 18216
rect 26620 18213 26648 18312
rect 28074 18300 28080 18312
rect 28132 18300 28138 18352
rect 29181 18343 29239 18349
rect 29181 18309 29193 18343
rect 29227 18340 29239 18343
rect 29362 18340 29368 18352
rect 29227 18312 29368 18340
rect 29227 18309 29239 18312
rect 29181 18303 29239 18309
rect 29362 18300 29368 18312
rect 29420 18300 29426 18352
rect 27341 18275 27399 18281
rect 27341 18241 27353 18275
rect 27387 18272 27399 18275
rect 27893 18275 27951 18281
rect 27893 18272 27905 18275
rect 27387 18244 27905 18272
rect 27387 18241 27399 18244
rect 27341 18235 27399 18241
rect 27893 18241 27905 18244
rect 27939 18241 27951 18275
rect 27893 18235 27951 18241
rect 27982 18232 27988 18284
rect 28040 18272 28046 18284
rect 28445 18275 28503 18281
rect 28445 18272 28457 18275
rect 28040 18244 28457 18272
rect 28040 18232 28046 18244
rect 28445 18241 28457 18244
rect 28491 18241 28503 18275
rect 28445 18235 28503 18241
rect 28718 18232 28724 18284
rect 28776 18272 28782 18284
rect 29641 18275 29699 18281
rect 29641 18272 29653 18275
rect 28776 18244 29653 18272
rect 28776 18232 28782 18244
rect 29641 18241 29653 18244
rect 29687 18241 29699 18275
rect 29641 18235 29699 18241
rect 26421 18207 26479 18213
rect 26421 18173 26433 18207
rect 26467 18173 26479 18207
rect 26421 18167 26479 18173
rect 26605 18207 26663 18213
rect 26605 18173 26617 18207
rect 26651 18173 26663 18207
rect 26605 18167 26663 18173
rect 27433 18207 27491 18213
rect 27433 18173 27445 18207
rect 27479 18173 27491 18207
rect 27433 18167 27491 18173
rect 27525 18207 27583 18213
rect 27525 18173 27537 18207
rect 27571 18204 27583 18207
rect 29730 18204 29736 18216
rect 27571 18176 29736 18204
rect 27571 18173 27583 18176
rect 27525 18167 27583 18173
rect 21634 18096 21640 18148
rect 21692 18136 21698 18148
rect 26436 18136 26464 18167
rect 27448 18136 27476 18167
rect 29730 18164 29736 18176
rect 29788 18164 29794 18216
rect 21692 18108 27476 18136
rect 29365 18139 29423 18145
rect 21692 18096 21698 18108
rect 29365 18105 29377 18139
rect 29411 18136 29423 18139
rect 29546 18136 29552 18148
rect 29411 18108 29552 18136
rect 29411 18105 29423 18108
rect 29365 18099 29423 18105
rect 29546 18096 29552 18108
rect 29604 18096 29610 18148
rect 21453 18071 21511 18077
rect 21453 18037 21465 18071
rect 21499 18037 21511 18071
rect 21453 18031 21511 18037
rect 26418 18028 26424 18080
rect 26476 18068 26482 18080
rect 26973 18071 27031 18077
rect 26973 18068 26985 18071
rect 26476 18040 26985 18068
rect 26476 18028 26482 18040
rect 26973 18037 26985 18040
rect 27019 18037 27031 18071
rect 26973 18031 27031 18037
rect 29454 18028 29460 18080
rect 29512 18068 29518 18080
rect 29733 18071 29791 18077
rect 29733 18068 29745 18071
rect 29512 18040 29745 18068
rect 29512 18028 29518 18040
rect 29733 18037 29745 18040
rect 29779 18037 29791 18071
rect 29733 18031 29791 18037
rect 1104 17978 31832 18000
rect 1104 17926 4182 17978
rect 4234 17926 4246 17978
rect 4298 17926 4310 17978
rect 4362 17926 4374 17978
rect 4426 17926 4438 17978
rect 4490 17926 4502 17978
rect 4554 17926 10182 17978
rect 10234 17926 10246 17978
rect 10298 17926 10310 17978
rect 10362 17926 10374 17978
rect 10426 17926 10438 17978
rect 10490 17926 10502 17978
rect 10554 17926 16182 17978
rect 16234 17926 16246 17978
rect 16298 17926 16310 17978
rect 16362 17926 16374 17978
rect 16426 17926 16438 17978
rect 16490 17926 16502 17978
rect 16554 17926 22182 17978
rect 22234 17926 22246 17978
rect 22298 17926 22310 17978
rect 22362 17926 22374 17978
rect 22426 17926 22438 17978
rect 22490 17926 22502 17978
rect 22554 17926 28182 17978
rect 28234 17926 28246 17978
rect 28298 17926 28310 17978
rect 28362 17926 28374 17978
rect 28426 17926 28438 17978
rect 28490 17926 28502 17978
rect 28554 17926 31832 17978
rect 1104 17904 31832 17926
rect 8389 17867 8447 17873
rect 8389 17833 8401 17867
rect 8435 17864 8447 17867
rect 8846 17864 8852 17876
rect 8435 17836 8852 17864
rect 8435 17833 8447 17836
rect 8389 17827 8447 17833
rect 8846 17824 8852 17836
rect 8904 17864 8910 17876
rect 9214 17864 9220 17876
rect 8904 17836 9220 17864
rect 8904 17824 8910 17836
rect 9214 17824 9220 17836
rect 9272 17824 9278 17876
rect 12713 17867 12771 17873
rect 12713 17833 12725 17867
rect 12759 17864 12771 17867
rect 13262 17864 13268 17876
rect 12759 17836 13268 17864
rect 12759 17833 12771 17836
rect 12713 17827 12771 17833
rect 13262 17824 13268 17836
rect 13320 17824 13326 17876
rect 14274 17824 14280 17876
rect 14332 17824 14338 17876
rect 15378 17824 15384 17876
rect 15436 17864 15442 17876
rect 20993 17867 21051 17873
rect 15436 17836 16436 17864
rect 15436 17824 15442 17836
rect 5810 17756 5816 17808
rect 5868 17756 5874 17808
rect 15286 17756 15292 17808
rect 15344 17796 15350 17808
rect 16408 17805 16436 17836
rect 20993 17833 21005 17867
rect 21039 17864 21051 17867
rect 21174 17864 21180 17876
rect 21039 17836 21180 17864
rect 21039 17833 21051 17836
rect 20993 17827 21051 17833
rect 21174 17824 21180 17836
rect 21232 17824 21238 17876
rect 21266 17824 21272 17876
rect 21324 17824 21330 17876
rect 16301 17799 16359 17805
rect 16301 17796 16313 17799
rect 15344 17768 16313 17796
rect 15344 17756 15350 17768
rect 16301 17765 16313 17768
rect 16347 17765 16359 17799
rect 16301 17759 16359 17765
rect 16393 17799 16451 17805
rect 16393 17765 16405 17799
rect 16439 17765 16451 17799
rect 16393 17759 16451 17765
rect 19797 17799 19855 17805
rect 19797 17765 19809 17799
rect 19843 17796 19855 17799
rect 21284 17796 21312 17824
rect 19843 17768 21312 17796
rect 19843 17765 19855 17768
rect 19797 17759 19855 17765
rect 30190 17756 30196 17808
rect 30248 17796 30254 17808
rect 30653 17799 30711 17805
rect 30653 17796 30665 17799
rect 30248 17768 30665 17796
rect 30248 17756 30254 17768
rect 30653 17765 30665 17768
rect 30699 17765 30711 17799
rect 30653 17759 30711 17765
rect 5828 17728 5856 17756
rect 5828 17700 6224 17728
rect 6196 17669 6224 17700
rect 12618 17688 12624 17740
rect 12676 17728 12682 17740
rect 13265 17731 13323 17737
rect 13265 17728 13277 17731
rect 12676 17700 13277 17728
rect 12676 17688 12682 17700
rect 13265 17697 13277 17700
rect 13311 17697 13323 17731
rect 13265 17691 13323 17697
rect 13449 17731 13507 17737
rect 13449 17697 13461 17731
rect 13495 17728 13507 17731
rect 13495 17700 14780 17728
rect 13495 17697 13507 17700
rect 13449 17691 13507 17697
rect 5629 17663 5687 17669
rect 5629 17660 5641 17663
rect 4816 17632 5641 17660
rect 4816 17536 4844 17632
rect 5629 17629 5641 17632
rect 5675 17660 5687 17663
rect 5813 17663 5871 17669
rect 5813 17660 5825 17663
rect 5675 17632 5825 17660
rect 5675 17629 5687 17632
rect 5629 17623 5687 17629
rect 5813 17629 5825 17632
rect 5859 17629 5871 17663
rect 5813 17623 5871 17629
rect 6181 17663 6239 17669
rect 6181 17629 6193 17663
rect 6227 17629 6239 17663
rect 6181 17623 6239 17629
rect 6914 17620 6920 17672
rect 6972 17660 6978 17672
rect 7282 17669 7288 17672
rect 7009 17663 7067 17669
rect 7009 17660 7021 17663
rect 6972 17632 7021 17660
rect 6972 17620 6978 17632
rect 7009 17629 7021 17632
rect 7055 17629 7067 17663
rect 7276 17660 7288 17669
rect 7243 17632 7288 17660
rect 7009 17623 7067 17629
rect 7276 17623 7288 17632
rect 7282 17620 7288 17623
rect 7340 17620 7346 17672
rect 12158 17620 12164 17672
rect 12216 17620 12222 17672
rect 12434 17620 12440 17672
rect 12492 17620 12498 17672
rect 12526 17620 12532 17672
rect 12584 17620 12590 17672
rect 14093 17663 14151 17669
rect 14093 17660 14105 17663
rect 13924 17632 14105 17660
rect 5718 17552 5724 17604
rect 5776 17592 5782 17604
rect 5997 17595 6055 17601
rect 5997 17592 6009 17595
rect 5776 17564 6009 17592
rect 5776 17552 5782 17564
rect 5997 17561 6009 17564
rect 6043 17561 6055 17595
rect 5997 17555 6055 17561
rect 6086 17552 6092 17604
rect 6144 17552 6150 17604
rect 12342 17552 12348 17604
rect 12400 17552 12406 17604
rect 4798 17484 4804 17536
rect 4856 17484 4862 17536
rect 5077 17527 5135 17533
rect 5077 17493 5089 17527
rect 5123 17524 5135 17527
rect 5350 17524 5356 17536
rect 5123 17496 5356 17524
rect 5123 17493 5135 17496
rect 5077 17487 5135 17493
rect 5350 17484 5356 17496
rect 5408 17484 5414 17536
rect 6362 17484 6368 17536
rect 6420 17484 6426 17536
rect 13538 17484 13544 17536
rect 13596 17484 13602 17536
rect 13924 17533 13952 17632
rect 14093 17629 14105 17632
rect 14139 17629 14151 17663
rect 14093 17623 14151 17629
rect 13909 17527 13967 17533
rect 13909 17493 13921 17527
rect 13955 17493 13967 17527
rect 13909 17487 13967 17493
rect 13998 17484 14004 17536
rect 14056 17524 14062 17536
rect 14461 17527 14519 17533
rect 14461 17524 14473 17527
rect 14056 17496 14473 17524
rect 14056 17484 14062 17496
rect 14461 17493 14473 17496
rect 14507 17493 14519 17527
rect 14752 17524 14780 17700
rect 14918 17688 14924 17740
rect 14976 17728 14982 17740
rect 15013 17731 15071 17737
rect 15013 17728 15025 17731
rect 14976 17700 15025 17728
rect 14976 17688 14982 17700
rect 15013 17697 15025 17700
rect 15059 17697 15071 17731
rect 15013 17691 15071 17697
rect 15470 17688 15476 17740
rect 15528 17728 15534 17740
rect 19978 17728 19984 17740
rect 15528 17700 16068 17728
rect 15528 17688 15534 17700
rect 16040 17669 16068 17700
rect 16224 17700 19380 17728
rect 16224 17669 16252 17700
rect 19352 17672 19380 17700
rect 19444 17700 19984 17728
rect 15841 17663 15899 17669
rect 15841 17629 15853 17663
rect 15887 17629 15899 17663
rect 15841 17623 15899 17629
rect 16025 17663 16083 17669
rect 16025 17629 16037 17663
rect 16071 17629 16083 17663
rect 16025 17623 16083 17629
rect 16209 17663 16267 17669
rect 16209 17629 16221 17663
rect 16255 17629 16267 17663
rect 16209 17623 16267 17629
rect 14829 17595 14887 17601
rect 14829 17561 14841 17595
rect 14875 17592 14887 17595
rect 15289 17595 15347 17601
rect 15289 17592 15301 17595
rect 14875 17564 15301 17592
rect 14875 17561 14887 17564
rect 14829 17555 14887 17561
rect 15289 17561 15301 17564
rect 15335 17561 15347 17595
rect 15289 17555 15347 17561
rect 15856 17536 15884 17623
rect 16482 17620 16488 17672
rect 16540 17620 16546 17672
rect 19245 17663 19303 17669
rect 19245 17629 19257 17663
rect 19291 17629 19303 17663
rect 19245 17623 19303 17629
rect 18414 17552 18420 17604
rect 18472 17552 18478 17604
rect 19260 17592 19288 17623
rect 19334 17620 19340 17672
rect 19392 17620 19398 17672
rect 19444 17669 19472 17700
rect 19978 17688 19984 17700
rect 20036 17728 20042 17740
rect 26878 17728 26884 17740
rect 20036 17700 26884 17728
rect 20036 17688 20042 17700
rect 26878 17688 26884 17700
rect 26936 17688 26942 17740
rect 29362 17688 29368 17740
rect 29420 17688 29426 17740
rect 29730 17688 29736 17740
rect 29788 17688 29794 17740
rect 19429 17663 19487 17669
rect 19429 17629 19441 17663
rect 19475 17629 19487 17663
rect 19429 17623 19487 17629
rect 19518 17620 19524 17672
rect 19576 17620 19582 17672
rect 19613 17663 19671 17669
rect 19613 17629 19625 17663
rect 19659 17660 19671 17663
rect 19794 17660 19800 17672
rect 19659 17632 19800 17660
rect 19659 17629 19671 17632
rect 19613 17623 19671 17629
rect 19794 17620 19800 17632
rect 19852 17620 19858 17672
rect 20438 17620 20444 17672
rect 20496 17620 20502 17672
rect 20714 17620 20720 17672
rect 20772 17620 20778 17672
rect 20809 17663 20867 17669
rect 20809 17629 20821 17663
rect 20855 17660 20867 17663
rect 20898 17660 20904 17672
rect 20855 17632 20904 17660
rect 20855 17629 20867 17632
rect 20809 17623 20867 17629
rect 20898 17620 20904 17632
rect 20956 17620 20962 17672
rect 21542 17620 21548 17672
rect 21600 17620 21606 17672
rect 23934 17620 23940 17672
rect 23992 17660 23998 17672
rect 24397 17663 24455 17669
rect 24397 17660 24409 17663
rect 23992 17632 24409 17660
rect 23992 17620 23998 17632
rect 24397 17629 24409 17632
rect 24443 17629 24455 17663
rect 30837 17663 30895 17669
rect 30837 17660 30849 17663
rect 24397 17623 24455 17629
rect 30300 17632 30849 17660
rect 19260 17564 19380 17592
rect 19352 17536 19380 17564
rect 20346 17552 20352 17604
rect 20404 17552 20410 17604
rect 20625 17595 20683 17601
rect 20625 17561 20637 17595
rect 20671 17592 20683 17595
rect 21560 17592 21588 17620
rect 21726 17592 21732 17604
rect 20671 17564 21732 17592
rect 20671 17561 20683 17564
rect 20625 17555 20683 17561
rect 21726 17552 21732 17564
rect 21784 17552 21790 17604
rect 14921 17527 14979 17533
rect 14921 17524 14933 17527
rect 14752 17496 14933 17524
rect 14461 17487 14519 17493
rect 14921 17493 14933 17496
rect 14967 17524 14979 17527
rect 15010 17524 15016 17536
rect 14967 17496 15016 17524
rect 14967 17493 14979 17496
rect 14921 17487 14979 17493
rect 15010 17484 15016 17496
rect 15068 17484 15074 17536
rect 15838 17484 15844 17536
rect 15896 17484 15902 17536
rect 17129 17527 17187 17533
rect 17129 17493 17141 17527
rect 17175 17524 17187 17527
rect 17862 17524 17868 17536
rect 17175 17496 17868 17524
rect 17175 17493 17187 17496
rect 17129 17487 17187 17493
rect 17862 17484 17868 17496
rect 17920 17484 17926 17536
rect 19334 17484 19340 17536
rect 19392 17524 19398 17536
rect 20364 17524 20392 17552
rect 19392 17496 20392 17524
rect 19392 17484 19398 17496
rect 25038 17484 25044 17536
rect 25096 17484 25102 17536
rect 28718 17484 28724 17536
rect 28776 17484 28782 17536
rect 28810 17484 28816 17536
rect 28868 17524 28874 17536
rect 29825 17527 29883 17533
rect 29825 17524 29837 17527
rect 28868 17496 29837 17524
rect 28868 17484 28874 17496
rect 29825 17493 29837 17496
rect 29871 17493 29883 17527
rect 29825 17487 29883 17493
rect 29914 17484 29920 17536
rect 29972 17484 29978 17536
rect 30300 17533 30328 17632
rect 30837 17629 30849 17632
rect 30883 17629 30895 17663
rect 30837 17623 30895 17629
rect 30285 17527 30343 17533
rect 30285 17493 30297 17527
rect 30331 17493 30343 17527
rect 30285 17487 30343 17493
rect 1104 17434 31832 17456
rect 1104 17382 4922 17434
rect 4974 17382 4986 17434
rect 5038 17382 5050 17434
rect 5102 17382 5114 17434
rect 5166 17382 5178 17434
rect 5230 17382 5242 17434
rect 5294 17382 10922 17434
rect 10974 17382 10986 17434
rect 11038 17382 11050 17434
rect 11102 17382 11114 17434
rect 11166 17382 11178 17434
rect 11230 17382 11242 17434
rect 11294 17382 16922 17434
rect 16974 17382 16986 17434
rect 17038 17382 17050 17434
rect 17102 17382 17114 17434
rect 17166 17382 17178 17434
rect 17230 17382 17242 17434
rect 17294 17382 22922 17434
rect 22974 17382 22986 17434
rect 23038 17382 23050 17434
rect 23102 17382 23114 17434
rect 23166 17382 23178 17434
rect 23230 17382 23242 17434
rect 23294 17382 28922 17434
rect 28974 17382 28986 17434
rect 29038 17382 29050 17434
rect 29102 17382 29114 17434
rect 29166 17382 29178 17434
rect 29230 17382 29242 17434
rect 29294 17382 31832 17434
rect 1104 17360 31832 17382
rect 4798 17280 4804 17332
rect 4856 17280 4862 17332
rect 5261 17323 5319 17329
rect 5261 17289 5273 17323
rect 5307 17320 5319 17323
rect 5350 17320 5356 17332
rect 5307 17292 5356 17320
rect 5307 17289 5319 17292
rect 5261 17283 5319 17289
rect 5350 17280 5356 17292
rect 5408 17280 5414 17332
rect 6362 17280 6368 17332
rect 6420 17320 6426 17332
rect 13265 17323 13323 17329
rect 6420 17292 9076 17320
rect 6420 17280 6426 17292
rect 6816 17255 6874 17261
rect 3436 17224 4016 17252
rect 3436 17193 3464 17224
rect 3988 17196 4016 17224
rect 6816 17221 6828 17255
rect 6862 17252 6874 17255
rect 7006 17252 7012 17264
rect 6862 17224 7012 17252
rect 6862 17221 6874 17224
rect 6816 17215 6874 17221
rect 7006 17212 7012 17224
rect 7064 17212 7070 17264
rect 8846 17212 8852 17264
rect 8904 17212 8910 17264
rect 3421 17187 3479 17193
rect 3421 17153 3433 17187
rect 3467 17153 3479 17187
rect 3421 17147 3479 17153
rect 3510 17144 3516 17196
rect 3568 17184 3574 17196
rect 3677 17187 3735 17193
rect 3677 17184 3689 17187
rect 3568 17156 3689 17184
rect 3568 17144 3574 17156
rect 3677 17153 3689 17156
rect 3723 17153 3735 17187
rect 3677 17147 3735 17153
rect 3970 17144 3976 17196
rect 4028 17144 4034 17196
rect 8754 17144 8760 17196
rect 8812 17144 8818 17196
rect 9048 17193 9076 17292
rect 13265 17289 13277 17323
rect 13311 17289 13323 17323
rect 13265 17283 13323 17289
rect 13357 17323 13415 17329
rect 13357 17289 13369 17323
rect 13403 17320 13415 17323
rect 13538 17320 13544 17332
rect 13403 17292 13544 17320
rect 13403 17289 13415 17292
rect 13357 17283 13415 17289
rect 13280 17252 13308 17283
rect 13538 17280 13544 17292
rect 13596 17280 13602 17332
rect 15473 17323 15531 17329
rect 15473 17289 15485 17323
rect 15519 17320 15531 17323
rect 15838 17320 15844 17332
rect 15519 17292 15844 17320
rect 15519 17289 15531 17292
rect 15473 17283 15531 17289
rect 15838 17280 15844 17292
rect 15896 17320 15902 17332
rect 16301 17323 16359 17329
rect 15896 17292 16160 17320
rect 15896 17280 15902 17292
rect 14338 17255 14396 17261
rect 14338 17252 14350 17255
rect 13280 17224 14350 17252
rect 14338 17221 14350 17224
rect 14384 17221 14396 17255
rect 14338 17215 14396 17221
rect 15194 17212 15200 17264
rect 15252 17252 15258 17264
rect 15746 17252 15752 17264
rect 15252 17224 15752 17252
rect 15252 17212 15258 17224
rect 15746 17212 15752 17224
rect 15804 17252 15810 17264
rect 16132 17261 16160 17292
rect 16301 17289 16313 17323
rect 16347 17320 16359 17323
rect 16482 17320 16488 17332
rect 16347 17292 16488 17320
rect 16347 17289 16359 17292
rect 16301 17283 16359 17289
rect 16482 17280 16488 17292
rect 16540 17280 16546 17332
rect 19061 17323 19119 17329
rect 19061 17289 19073 17323
rect 19107 17320 19119 17323
rect 19334 17320 19340 17332
rect 19107 17292 19340 17320
rect 19107 17289 19119 17292
rect 19061 17283 19119 17289
rect 19334 17280 19340 17292
rect 19392 17280 19398 17332
rect 24857 17323 24915 17329
rect 24857 17289 24869 17323
rect 24903 17320 24915 17323
rect 25038 17320 25044 17332
rect 24903 17292 25044 17320
rect 24903 17289 24915 17292
rect 24857 17283 24915 17289
rect 25038 17280 25044 17292
rect 25096 17280 25102 17332
rect 26234 17280 26240 17332
rect 26292 17320 26298 17332
rect 27154 17320 27160 17332
rect 26292 17292 27160 17320
rect 26292 17280 26298 17292
rect 27154 17280 27160 17292
rect 27212 17280 27218 17332
rect 28445 17323 28503 17329
rect 28445 17289 28457 17323
rect 28491 17320 28503 17323
rect 28718 17320 28724 17332
rect 28491 17292 28724 17320
rect 28491 17289 28503 17292
rect 28445 17283 28503 17289
rect 28718 17280 28724 17292
rect 28776 17280 28782 17332
rect 28810 17280 28816 17332
rect 28868 17280 28874 17332
rect 28905 17323 28963 17329
rect 28905 17289 28917 17323
rect 28951 17320 28963 17323
rect 29178 17320 29184 17332
rect 28951 17292 29184 17320
rect 28951 17289 28963 17292
rect 28905 17283 28963 17289
rect 29178 17280 29184 17292
rect 29236 17320 29242 17332
rect 29362 17320 29368 17332
rect 29236 17292 29368 17320
rect 29236 17280 29242 17292
rect 29362 17280 29368 17292
rect 29420 17280 29426 17332
rect 29914 17280 29920 17332
rect 29972 17320 29978 17332
rect 30377 17323 30435 17329
rect 30377 17320 30389 17323
rect 29972 17292 30389 17320
rect 29972 17280 29978 17292
rect 30377 17289 30389 17292
rect 30423 17289 30435 17323
rect 30377 17283 30435 17289
rect 31113 17323 31171 17329
rect 31113 17289 31125 17323
rect 31159 17289 31171 17323
rect 31113 17283 31171 17289
rect 15933 17255 15991 17261
rect 15933 17252 15945 17255
rect 15804 17224 15945 17252
rect 15804 17212 15810 17224
rect 15933 17221 15945 17224
rect 15979 17221 15991 17255
rect 15933 17215 15991 17221
rect 16117 17255 16175 17261
rect 16117 17221 16129 17255
rect 16163 17221 16175 17255
rect 16117 17215 16175 17221
rect 19794 17212 19800 17264
rect 19852 17252 19858 17264
rect 20346 17252 20352 17264
rect 19852 17224 20352 17252
rect 19852 17212 19858 17224
rect 20346 17212 20352 17224
rect 20404 17252 20410 17264
rect 20404 17224 23796 17252
rect 20404 17212 20410 17224
rect 9033 17187 9091 17193
rect 9033 17153 9045 17187
rect 9079 17153 9091 17187
rect 9033 17147 9091 17153
rect 10413 17187 10471 17193
rect 10413 17153 10425 17187
rect 10459 17184 10471 17187
rect 10594 17184 10600 17196
rect 10459 17156 10600 17184
rect 10459 17153 10471 17156
rect 10413 17147 10471 17153
rect 10594 17144 10600 17156
rect 10652 17144 10658 17196
rect 13081 17187 13139 17193
rect 13081 17153 13093 17187
rect 13127 17184 13139 17187
rect 13998 17184 14004 17196
rect 13127 17156 14004 17184
rect 13127 17153 13139 17156
rect 13081 17147 13139 17153
rect 13998 17144 14004 17156
rect 14056 17144 14062 17196
rect 14093 17187 14151 17193
rect 14093 17153 14105 17187
rect 14139 17184 14151 17187
rect 14182 17184 14188 17196
rect 14139 17156 14188 17184
rect 14139 17153 14151 17156
rect 14093 17147 14151 17153
rect 14182 17144 14188 17156
rect 14240 17144 14246 17196
rect 17310 17144 17316 17196
rect 17368 17184 17374 17196
rect 17681 17187 17739 17193
rect 17681 17184 17693 17187
rect 17368 17156 17693 17184
rect 17368 17144 17374 17156
rect 17681 17153 17693 17156
rect 17727 17153 17739 17187
rect 17681 17147 17739 17153
rect 17948 17187 18006 17193
rect 17948 17153 17960 17187
rect 17994 17184 18006 17187
rect 18230 17184 18236 17196
rect 17994 17156 18236 17184
rect 17994 17153 18006 17156
rect 17948 17147 18006 17153
rect 18230 17144 18236 17156
rect 18288 17144 18294 17196
rect 22465 17187 22523 17193
rect 22465 17153 22477 17187
rect 22511 17184 22523 17187
rect 22646 17184 22652 17196
rect 22511 17156 22652 17184
rect 22511 17153 22523 17156
rect 22465 17147 22523 17153
rect 22646 17144 22652 17156
rect 22704 17144 22710 17196
rect 4614 17076 4620 17128
rect 4672 17076 4678 17128
rect 5350 17076 5356 17128
rect 5408 17076 5414 17128
rect 5445 17119 5503 17125
rect 5445 17085 5457 17119
rect 5491 17085 5503 17119
rect 5445 17079 5503 17085
rect 6549 17119 6607 17125
rect 6549 17085 6561 17119
rect 6595 17085 6607 17119
rect 6549 17079 6607 17085
rect 8665 17119 8723 17125
rect 8665 17085 8677 17119
rect 8711 17116 8723 17119
rect 8711 17088 9076 17116
rect 8711 17085 8723 17088
rect 8665 17079 8723 17085
rect 4632 17048 4660 17076
rect 5460 17048 5488 17079
rect 4632 17020 5488 17048
rect 4890 16940 4896 16992
rect 4948 16940 4954 16992
rect 6564 16980 6592 17079
rect 7929 17051 7987 17057
rect 7929 17017 7941 17051
rect 7975 17048 7987 17051
rect 8680 17048 8708 17079
rect 7975 17020 8708 17048
rect 7975 17017 7987 17020
rect 7929 17011 7987 17017
rect 9048 16992 9076 17088
rect 13906 17076 13912 17128
rect 13964 17076 13970 17128
rect 23566 17076 23572 17128
rect 23624 17076 23630 17128
rect 23768 17116 23796 17224
rect 23952 17224 26648 17252
rect 23952 17196 23980 17224
rect 23842 17144 23848 17196
rect 23900 17144 23906 17196
rect 23934 17144 23940 17196
rect 23992 17144 23998 17196
rect 24765 17187 24823 17193
rect 24044 17156 24716 17184
rect 24044 17116 24072 17156
rect 23768 17088 24072 17116
rect 24581 17119 24639 17125
rect 24581 17085 24593 17119
rect 24627 17085 24639 17119
rect 24688 17116 24716 17156
rect 24765 17153 24777 17187
rect 24811 17184 24823 17187
rect 26050 17184 26056 17196
rect 24811 17156 26056 17184
rect 24811 17153 24823 17156
rect 24765 17147 24823 17153
rect 26050 17144 26056 17156
rect 26108 17144 26114 17196
rect 26234 17144 26240 17196
rect 26292 17144 26298 17196
rect 26620 17193 26648 17224
rect 26878 17212 26884 17264
rect 26936 17212 26942 17264
rect 27614 17212 27620 17264
rect 27672 17252 27678 17264
rect 28353 17255 28411 17261
rect 28353 17252 28365 17255
rect 27672 17224 28365 17252
rect 27672 17212 27678 17224
rect 28353 17221 28365 17224
rect 28399 17252 28411 17255
rect 28828 17252 28856 17280
rect 28399 17224 28856 17252
rect 28399 17221 28411 17224
rect 28353 17215 28411 17221
rect 29086 17212 29092 17264
rect 29144 17252 29150 17264
rect 29454 17252 29460 17264
rect 29144 17224 29460 17252
rect 29144 17212 29150 17224
rect 29454 17212 29460 17224
rect 29512 17212 29518 17264
rect 29822 17252 29828 17264
rect 29656 17224 29828 17252
rect 26329 17187 26387 17193
rect 26329 17153 26341 17187
rect 26375 17153 26387 17187
rect 26329 17147 26387 17153
rect 26421 17187 26479 17193
rect 26421 17153 26433 17187
rect 26467 17153 26479 17187
rect 26421 17147 26479 17153
rect 26605 17187 26663 17193
rect 26605 17153 26617 17187
rect 26651 17153 26663 17187
rect 26605 17147 26663 17153
rect 24688 17088 25820 17116
rect 24581 17079 24639 17085
rect 9122 17008 9128 17060
rect 9180 17048 9186 17060
rect 9180 17020 12112 17048
rect 9180 17008 9186 17020
rect 12084 16992 12112 17020
rect 19886 17008 19892 17060
rect 19944 17048 19950 17060
rect 20254 17048 20260 17060
rect 19944 17020 20260 17048
rect 19944 17008 19950 17020
rect 20254 17008 20260 17020
rect 20312 17048 20318 17060
rect 24596 17048 24624 17079
rect 20312 17020 24624 17048
rect 25225 17051 25283 17057
rect 20312 17008 20318 17020
rect 25225 17017 25237 17051
rect 25271 17048 25283 17051
rect 25682 17048 25688 17060
rect 25271 17020 25688 17048
rect 25271 17017 25283 17020
rect 25225 17011 25283 17017
rect 25682 17008 25688 17020
rect 25740 17008 25746 17060
rect 25792 17048 25820 17088
rect 25866 17076 25872 17128
rect 25924 17116 25930 17128
rect 26344 17116 26372 17147
rect 25924 17088 26372 17116
rect 26436 17116 26464 17147
rect 26896 17116 26924 17212
rect 29656 17196 29684 17224
rect 29822 17212 29828 17224
rect 29880 17212 29886 17264
rect 30040 17255 30098 17261
rect 30040 17221 30052 17255
rect 30086 17252 30098 17255
rect 31128 17252 31156 17283
rect 30086 17224 31156 17252
rect 30086 17221 30098 17224
rect 30040 17215 30098 17221
rect 28074 17144 28080 17196
rect 28132 17184 28138 17196
rect 29638 17184 29644 17196
rect 28132 17156 29644 17184
rect 28132 17144 28138 17156
rect 28276 17125 28304 17156
rect 29638 17144 29644 17156
rect 29696 17144 29702 17196
rect 30285 17187 30343 17193
rect 30285 17153 30297 17187
rect 30331 17184 30343 17187
rect 30558 17184 30564 17196
rect 30331 17156 30564 17184
rect 30331 17153 30343 17156
rect 30285 17147 30343 17153
rect 30558 17144 30564 17156
rect 30616 17144 30622 17196
rect 31297 17187 31355 17193
rect 31297 17184 31309 17187
rect 30668 17156 31309 17184
rect 26436 17088 26924 17116
rect 28261 17119 28319 17125
rect 25924 17076 25930 17088
rect 28261 17085 28273 17119
rect 28307 17085 28319 17119
rect 28261 17079 28319 17085
rect 26234 17048 26240 17060
rect 25792 17020 26240 17048
rect 26234 17008 26240 17020
rect 26292 17008 26298 17060
rect 6914 16980 6920 16992
rect 6564 16952 6920 16980
rect 6914 16940 6920 16952
rect 6972 16980 6978 16992
rect 7834 16980 7840 16992
rect 6972 16952 7840 16980
rect 6972 16940 6978 16952
rect 7834 16940 7840 16952
rect 7892 16940 7898 16992
rect 8018 16940 8024 16992
rect 8076 16940 8082 16992
rect 9030 16940 9036 16992
rect 9088 16940 9094 16992
rect 9217 16983 9275 16989
rect 9217 16949 9229 16983
rect 9263 16980 9275 16983
rect 9674 16980 9680 16992
rect 9263 16952 9680 16980
rect 9263 16949 9275 16952
rect 9217 16943 9275 16949
rect 9674 16940 9680 16952
rect 9732 16940 9738 16992
rect 10042 16940 10048 16992
rect 10100 16980 10106 16992
rect 10229 16983 10287 16989
rect 10229 16980 10241 16983
rect 10100 16952 10241 16980
rect 10100 16940 10106 16952
rect 10229 16949 10241 16952
rect 10275 16949 10287 16983
rect 10229 16943 10287 16949
rect 12066 16940 12072 16992
rect 12124 16940 12130 16992
rect 22094 16940 22100 16992
rect 22152 16980 22158 16992
rect 22281 16983 22339 16989
rect 22281 16980 22293 16983
rect 22152 16952 22293 16980
rect 22152 16940 22158 16952
rect 22281 16949 22293 16952
rect 22327 16949 22339 16983
rect 22281 16943 22339 16949
rect 22738 16940 22744 16992
rect 22796 16980 22802 16992
rect 22925 16983 22983 16989
rect 22925 16980 22937 16983
rect 22796 16952 22937 16980
rect 22796 16940 22802 16952
rect 22925 16949 22937 16952
rect 22971 16949 22983 16983
rect 22925 16943 22983 16949
rect 24026 16940 24032 16992
rect 24084 16940 24090 16992
rect 25314 16940 25320 16992
rect 25372 16940 25378 16992
rect 25774 16940 25780 16992
rect 25832 16980 25838 16992
rect 26053 16983 26111 16989
rect 26053 16980 26065 16983
rect 25832 16952 26065 16980
rect 25832 16940 25838 16952
rect 26053 16949 26065 16952
rect 26099 16949 26111 16983
rect 26053 16943 26111 16949
rect 28813 16983 28871 16989
rect 28813 16949 28825 16983
rect 28859 16980 28871 16983
rect 30668 16980 30696 17156
rect 31297 17153 31309 17156
rect 31343 17153 31355 17187
rect 31297 17147 31355 17153
rect 30926 17076 30932 17128
rect 30984 17076 30990 17128
rect 28859 16952 30696 16980
rect 28859 16949 28871 16952
rect 28813 16943 28871 16949
rect 1104 16890 31832 16912
rect 1104 16838 4182 16890
rect 4234 16838 4246 16890
rect 4298 16838 4310 16890
rect 4362 16838 4374 16890
rect 4426 16838 4438 16890
rect 4490 16838 4502 16890
rect 4554 16838 10182 16890
rect 10234 16838 10246 16890
rect 10298 16838 10310 16890
rect 10362 16838 10374 16890
rect 10426 16838 10438 16890
rect 10490 16838 10502 16890
rect 10554 16838 16182 16890
rect 16234 16838 16246 16890
rect 16298 16838 16310 16890
rect 16362 16838 16374 16890
rect 16426 16838 16438 16890
rect 16490 16838 16502 16890
rect 16554 16838 22182 16890
rect 22234 16838 22246 16890
rect 22298 16838 22310 16890
rect 22362 16838 22374 16890
rect 22426 16838 22438 16890
rect 22490 16838 22502 16890
rect 22554 16838 28182 16890
rect 28234 16838 28246 16890
rect 28298 16838 28310 16890
rect 28362 16838 28374 16890
rect 28426 16838 28438 16890
rect 28490 16838 28502 16890
rect 28554 16838 31832 16890
rect 1104 16816 31832 16838
rect 3329 16779 3387 16785
rect 3329 16745 3341 16779
rect 3375 16776 3387 16779
rect 3510 16776 3516 16788
rect 3375 16748 3516 16776
rect 3375 16745 3387 16748
rect 3329 16739 3387 16745
rect 3510 16736 3516 16748
rect 3568 16736 3574 16788
rect 3970 16776 3976 16788
rect 3804 16748 3976 16776
rect 3804 16649 3832 16748
rect 3970 16736 3976 16748
rect 4028 16736 4034 16788
rect 6917 16779 6975 16785
rect 6917 16745 6929 16779
rect 6963 16776 6975 16779
rect 7006 16776 7012 16788
rect 6963 16748 7012 16776
rect 6963 16745 6975 16748
rect 6917 16739 6975 16745
rect 7006 16736 7012 16748
rect 7064 16736 7070 16788
rect 8754 16736 8760 16788
rect 8812 16776 8818 16788
rect 8812 16748 12020 16776
rect 8812 16736 8818 16748
rect 5350 16668 5356 16720
rect 5408 16708 5414 16720
rect 9122 16708 9128 16720
rect 5408 16680 6868 16708
rect 5408 16668 5414 16680
rect 3789 16643 3847 16649
rect 3789 16609 3801 16643
rect 3835 16609 3847 16643
rect 3789 16603 3847 16609
rect 5905 16643 5963 16649
rect 5905 16609 5917 16643
rect 5951 16640 5963 16643
rect 6086 16640 6092 16652
rect 5951 16612 6092 16640
rect 5951 16609 5963 16612
rect 5905 16603 5963 16609
rect 3145 16575 3203 16581
rect 3145 16541 3157 16575
rect 3191 16541 3203 16575
rect 3145 16535 3203 16541
rect 3160 16504 3188 16535
rect 3418 16532 3424 16584
rect 3476 16532 3482 16584
rect 4890 16572 4896 16584
rect 3528 16544 4896 16572
rect 3528 16504 3556 16544
rect 4890 16532 4896 16544
rect 4948 16532 4954 16584
rect 4034 16507 4092 16513
rect 4034 16504 4046 16507
rect 3160 16476 3556 16504
rect 3620 16476 4046 16504
rect 3620 16445 3648 16476
rect 4034 16473 4046 16476
rect 4080 16473 4092 16507
rect 4034 16467 4092 16473
rect 4614 16464 4620 16516
rect 4672 16504 4678 16516
rect 5261 16507 5319 16513
rect 5261 16504 5273 16507
rect 4672 16476 5273 16504
rect 4672 16464 4678 16476
rect 5261 16473 5273 16476
rect 5307 16473 5319 16507
rect 5261 16467 5319 16473
rect 3605 16439 3663 16445
rect 3605 16405 3617 16439
rect 3651 16405 3663 16439
rect 3605 16399 3663 16405
rect 5169 16439 5227 16445
rect 5169 16405 5181 16439
rect 5215 16436 5227 16439
rect 5920 16436 5948 16603
rect 6086 16600 6092 16612
rect 6144 16600 6150 16652
rect 6840 16640 6868 16680
rect 7300 16680 9128 16708
rect 7300 16640 7328 16680
rect 9122 16668 9128 16680
rect 9180 16668 9186 16720
rect 11149 16711 11207 16717
rect 11149 16677 11161 16711
rect 11195 16708 11207 16711
rect 11698 16708 11704 16720
rect 11195 16680 11704 16708
rect 11195 16677 11207 16680
rect 11149 16671 11207 16677
rect 11698 16668 11704 16680
rect 11756 16708 11762 16720
rect 11992 16708 12020 16748
rect 12066 16736 12072 16788
rect 12124 16776 12130 16788
rect 13078 16776 13084 16788
rect 12124 16748 13084 16776
rect 12124 16736 12130 16748
rect 13078 16736 13084 16748
rect 13136 16776 13142 16788
rect 15194 16776 15200 16788
rect 13136 16748 15200 16776
rect 13136 16736 13142 16748
rect 15194 16736 15200 16748
rect 15252 16736 15258 16788
rect 18230 16736 18236 16788
rect 18288 16736 18294 16788
rect 19150 16736 19156 16788
rect 19208 16776 19214 16788
rect 19208 16748 23612 16776
rect 19208 16736 19214 16748
rect 14642 16708 14648 16720
rect 11756 16680 11836 16708
rect 11992 16680 14648 16708
rect 11756 16668 11762 16680
rect 6840 16612 7328 16640
rect 6840 16584 6868 16612
rect 6822 16532 6828 16584
rect 6880 16532 6886 16584
rect 7101 16575 7159 16581
rect 7101 16541 7113 16575
rect 7147 16572 7159 16575
rect 7147 16544 7236 16572
rect 7147 16541 7159 16544
rect 7101 16535 7159 16541
rect 7208 16445 7236 16544
rect 7300 16504 7328 16612
rect 7374 16600 7380 16652
rect 7432 16640 7438 16652
rect 7745 16643 7803 16649
rect 7745 16640 7757 16643
rect 7432 16612 7757 16640
rect 7432 16600 7438 16612
rect 7745 16609 7757 16612
rect 7791 16609 7803 16643
rect 7745 16603 7803 16609
rect 7834 16600 7840 16652
rect 7892 16640 7898 16652
rect 11808 16649 11836 16680
rect 14642 16668 14648 16680
rect 14700 16668 14706 16720
rect 9769 16643 9827 16649
rect 9769 16640 9781 16643
rect 7892 16612 9781 16640
rect 7892 16600 7898 16612
rect 9769 16609 9781 16612
rect 9815 16609 9827 16643
rect 9769 16603 9827 16609
rect 11793 16643 11851 16649
rect 11793 16609 11805 16643
rect 11839 16609 11851 16643
rect 11793 16603 11851 16609
rect 14182 16600 14188 16652
rect 14240 16640 14246 16652
rect 14366 16640 14372 16652
rect 14240 16612 14372 16640
rect 14240 16600 14246 16612
rect 14366 16600 14372 16612
rect 14424 16600 14430 16652
rect 23584 16649 23612 16748
rect 23842 16736 23848 16788
rect 23900 16776 23906 16788
rect 24213 16779 24271 16785
rect 24213 16776 24225 16779
rect 23900 16748 24225 16776
rect 23900 16736 23906 16748
rect 24213 16745 24225 16748
rect 24259 16745 24271 16779
rect 24213 16739 24271 16745
rect 25777 16779 25835 16785
rect 25777 16745 25789 16779
rect 25823 16776 25835 16779
rect 25866 16776 25872 16788
rect 25823 16748 25872 16776
rect 25823 16745 25835 16748
rect 25777 16739 25835 16745
rect 25866 16736 25872 16748
rect 25924 16736 25930 16788
rect 28626 16736 28632 16788
rect 28684 16776 28690 16788
rect 28684 16748 28994 16776
rect 28684 16736 28690 16748
rect 27154 16668 27160 16720
rect 27212 16708 27218 16720
rect 28721 16711 28779 16717
rect 28721 16708 28733 16711
rect 27212 16680 28733 16708
rect 27212 16668 27218 16680
rect 28721 16677 28733 16680
rect 28767 16677 28779 16711
rect 28966 16708 28994 16748
rect 29454 16736 29460 16788
rect 29512 16776 29518 16788
rect 29914 16776 29920 16788
rect 29512 16748 29920 16776
rect 29512 16736 29518 16748
rect 29914 16736 29920 16748
rect 29972 16736 29978 16788
rect 28966 16680 29592 16708
rect 28721 16671 28779 16677
rect 23569 16643 23627 16649
rect 23569 16609 23581 16643
rect 23615 16609 23627 16643
rect 23569 16603 23627 16609
rect 24397 16643 24455 16649
rect 24397 16609 24409 16643
rect 24443 16640 24455 16643
rect 24443 16612 24532 16640
rect 24443 16609 24455 16612
rect 24397 16603 24455 16609
rect 7561 16575 7619 16581
rect 7561 16541 7573 16575
rect 7607 16572 7619 16575
rect 8018 16572 8024 16584
rect 7607 16544 8024 16572
rect 7607 16541 7619 16544
rect 7561 16535 7619 16541
rect 8018 16532 8024 16544
rect 8076 16532 8082 16584
rect 10042 16581 10048 16584
rect 10036 16572 10048 16581
rect 10003 16544 10048 16572
rect 10036 16535 10048 16544
rect 10042 16532 10048 16535
rect 10100 16532 10106 16584
rect 7653 16507 7711 16513
rect 7653 16504 7665 16507
rect 7300 16476 7665 16504
rect 7653 16473 7665 16476
rect 7699 16473 7711 16507
rect 14200 16504 14228 16600
rect 18417 16575 18475 16581
rect 18417 16541 18429 16575
rect 18463 16572 18475 16575
rect 18966 16572 18972 16584
rect 18463 16544 18972 16572
rect 18463 16541 18475 16544
rect 18417 16535 18475 16541
rect 18966 16532 18972 16544
rect 19024 16532 19030 16584
rect 21542 16532 21548 16584
rect 21600 16572 21606 16584
rect 22094 16581 22100 16584
rect 21821 16575 21879 16581
rect 21821 16572 21833 16575
rect 21600 16544 21833 16572
rect 21600 16532 21606 16544
rect 21821 16541 21833 16544
rect 21867 16541 21879 16575
rect 21821 16535 21879 16541
rect 22088 16535 22100 16581
rect 22152 16572 22158 16584
rect 23753 16575 23811 16581
rect 22152 16544 22188 16572
rect 22094 16532 22100 16535
rect 22152 16532 22158 16544
rect 23753 16541 23765 16575
rect 23799 16572 23811 16575
rect 23842 16572 23848 16584
rect 23799 16544 23848 16572
rect 23799 16541 23811 16544
rect 23753 16535 23811 16541
rect 23842 16532 23848 16544
rect 23900 16532 23906 16584
rect 24026 16532 24032 16584
rect 24084 16532 24090 16584
rect 24504 16572 24532 16612
rect 29086 16600 29092 16652
rect 29144 16600 29150 16652
rect 29178 16600 29184 16652
rect 29236 16640 29242 16652
rect 29564 16649 29592 16680
rect 29549 16643 29607 16649
rect 29236 16612 29315 16640
rect 29236 16600 29242 16612
rect 25590 16572 25596 16584
rect 24504 16544 25596 16572
rect 25590 16532 25596 16544
rect 25648 16532 25654 16584
rect 25682 16532 25688 16584
rect 25740 16572 25746 16584
rect 28902 16581 28908 16584
rect 26053 16575 26111 16581
rect 26053 16572 26065 16575
rect 25740 16544 26065 16572
rect 25740 16532 25746 16544
rect 26053 16541 26065 16544
rect 26099 16541 26111 16575
rect 28900 16572 28908 16581
rect 28863 16544 28908 16572
rect 26053 16535 26111 16541
rect 28900 16535 28908 16544
rect 28902 16532 28908 16535
rect 28960 16532 28966 16584
rect 28997 16575 29055 16581
rect 28997 16541 29009 16575
rect 29043 16572 29055 16575
rect 29104 16572 29132 16600
rect 29287 16581 29315 16612
rect 29549 16609 29561 16643
rect 29595 16609 29607 16643
rect 29549 16603 29607 16609
rect 29043 16544 29132 16572
rect 29272 16575 29330 16581
rect 29043 16541 29055 16544
rect 28997 16535 29055 16541
rect 29272 16541 29284 16575
rect 29318 16541 29330 16575
rect 29272 16535 29330 16541
rect 29365 16575 29423 16581
rect 29365 16541 29377 16575
rect 29411 16572 29423 16575
rect 29454 16572 29460 16584
rect 29411 16544 29460 16572
rect 29411 16541 29423 16544
rect 29365 16535 29423 16541
rect 29454 16532 29460 16544
rect 29512 16532 29518 16584
rect 29816 16575 29874 16581
rect 29816 16541 29828 16575
rect 29862 16572 29874 16575
rect 30190 16572 30196 16584
rect 29862 16544 30196 16572
rect 29862 16541 29874 16544
rect 29816 16535 29874 16541
rect 30190 16532 30196 16544
rect 30248 16532 30254 16584
rect 30926 16532 30932 16584
rect 30984 16532 30990 16584
rect 7653 16467 7711 16473
rect 9600 16476 14228 16504
rect 24044 16504 24072 16532
rect 24642 16507 24700 16513
rect 24642 16504 24654 16507
rect 24044 16476 24654 16504
rect 9600 16448 9628 16476
rect 24642 16473 24654 16476
rect 24688 16473 24700 16507
rect 24642 16467 24700 16473
rect 25314 16464 25320 16516
rect 25372 16464 25378 16516
rect 29089 16507 29147 16513
rect 29089 16473 29101 16507
rect 29135 16504 29147 16507
rect 30650 16504 30656 16516
rect 29135 16476 30656 16504
rect 29135 16473 29147 16476
rect 29089 16467 29147 16473
rect 30650 16464 30656 16476
rect 30708 16464 30714 16516
rect 5215 16408 5948 16436
rect 7193 16439 7251 16445
rect 5215 16405 5227 16408
rect 5169 16399 5227 16405
rect 7193 16405 7205 16439
rect 7239 16405 7251 16439
rect 7193 16399 7251 16405
rect 9582 16396 9588 16448
rect 9640 16396 9646 16448
rect 11241 16439 11299 16445
rect 11241 16405 11253 16439
rect 11287 16436 11299 16439
rect 11330 16436 11336 16448
rect 11287 16408 11336 16436
rect 11287 16405 11299 16408
rect 11241 16399 11299 16405
rect 11330 16396 11336 16408
rect 11388 16396 11394 16448
rect 23201 16439 23259 16445
rect 23201 16405 23213 16439
rect 23247 16436 23259 16439
rect 23382 16436 23388 16448
rect 23247 16408 23388 16436
rect 23247 16405 23259 16408
rect 23201 16399 23259 16405
rect 23382 16396 23388 16408
rect 23440 16396 23446 16448
rect 23845 16439 23903 16445
rect 23845 16405 23857 16439
rect 23891 16436 23903 16439
rect 25332 16436 25360 16464
rect 23891 16408 25360 16436
rect 23891 16405 23903 16408
rect 23845 16399 23903 16405
rect 25866 16396 25872 16448
rect 25924 16396 25930 16448
rect 30944 16445 30972 16532
rect 30929 16439 30987 16445
rect 30929 16405 30941 16439
rect 30975 16405 30987 16439
rect 30929 16399 30987 16405
rect 1104 16346 31832 16368
rect 1104 16294 4922 16346
rect 4974 16294 4986 16346
rect 5038 16294 5050 16346
rect 5102 16294 5114 16346
rect 5166 16294 5178 16346
rect 5230 16294 5242 16346
rect 5294 16294 10922 16346
rect 10974 16294 10986 16346
rect 11038 16294 11050 16346
rect 11102 16294 11114 16346
rect 11166 16294 11178 16346
rect 11230 16294 11242 16346
rect 11294 16294 16922 16346
rect 16974 16294 16986 16346
rect 17038 16294 17050 16346
rect 17102 16294 17114 16346
rect 17166 16294 17178 16346
rect 17230 16294 17242 16346
rect 17294 16294 22922 16346
rect 22974 16294 22986 16346
rect 23038 16294 23050 16346
rect 23102 16294 23114 16346
rect 23166 16294 23178 16346
rect 23230 16294 23242 16346
rect 23294 16294 28922 16346
rect 28974 16294 28986 16346
rect 29038 16294 29050 16346
rect 29102 16294 29114 16346
rect 29166 16294 29178 16346
rect 29230 16294 29242 16346
rect 29294 16294 31832 16346
rect 1104 16272 31832 16294
rect 3418 16192 3424 16244
rect 3476 16232 3482 16244
rect 4249 16235 4307 16241
rect 4249 16232 4261 16235
rect 3476 16204 4261 16232
rect 3476 16192 3482 16204
rect 4249 16201 4261 16204
rect 4295 16201 4307 16235
rect 4249 16195 4307 16201
rect 4614 16192 4620 16244
rect 4672 16192 4678 16244
rect 4709 16235 4767 16241
rect 4709 16201 4721 16235
rect 4755 16232 4767 16235
rect 5350 16232 5356 16244
rect 4755 16204 5356 16232
rect 4755 16201 4767 16204
rect 4709 16195 4767 16201
rect 5350 16192 5356 16204
rect 5408 16192 5414 16244
rect 9490 16232 9496 16244
rect 9232 16204 9496 16232
rect 9232 16173 9260 16204
rect 9490 16192 9496 16204
rect 9548 16192 9554 16244
rect 10505 16235 10563 16241
rect 10505 16201 10517 16235
rect 10551 16232 10563 16235
rect 10594 16232 10600 16244
rect 10551 16204 10600 16232
rect 10551 16201 10563 16204
rect 10505 16195 10563 16201
rect 10594 16192 10600 16204
rect 10652 16192 10658 16244
rect 10873 16235 10931 16241
rect 10873 16201 10885 16235
rect 10919 16232 10931 16235
rect 11330 16232 11336 16244
rect 10919 16204 11336 16232
rect 10919 16201 10931 16204
rect 10873 16195 10931 16201
rect 11330 16192 11336 16204
rect 11388 16192 11394 16244
rect 21637 16235 21695 16241
rect 11624 16204 21588 16232
rect 9217 16167 9275 16173
rect 9217 16133 9229 16167
rect 9263 16133 9275 16167
rect 11517 16167 11575 16173
rect 11517 16164 11529 16167
rect 9217 16127 9275 16133
rect 9968 16136 11529 16164
rect 8938 16056 8944 16108
rect 8996 16056 9002 16108
rect 9030 16056 9036 16108
rect 9088 16056 9094 16108
rect 9306 16056 9312 16108
rect 9364 16056 9370 16108
rect 9447 16099 9505 16105
rect 9447 16065 9459 16099
rect 9493 16096 9505 16099
rect 9582 16096 9588 16108
rect 9493 16068 9588 16096
rect 9493 16065 9505 16068
rect 9447 16059 9505 16065
rect 9582 16056 9588 16068
rect 9640 16056 9646 16108
rect 9674 16056 9680 16108
rect 9732 16056 9738 16108
rect 9968 16105 9996 16136
rect 11517 16133 11529 16136
rect 11563 16133 11575 16167
rect 11517 16127 11575 16133
rect 9953 16099 10011 16105
rect 9953 16065 9965 16099
rect 9999 16065 10011 16099
rect 9953 16059 10011 16065
rect 10229 16099 10287 16105
rect 10229 16065 10241 16099
rect 10275 16096 10287 16099
rect 11624 16096 11652 16204
rect 11698 16124 11704 16176
rect 11756 16124 11762 16176
rect 12406 16136 15792 16164
rect 10275 16068 11652 16096
rect 10275 16065 10287 16068
rect 10229 16059 10287 16065
rect 11790 16056 11796 16108
rect 11848 16096 11854 16108
rect 11885 16099 11943 16105
rect 11885 16096 11897 16099
rect 11848 16068 11897 16096
rect 11848 16056 11854 16068
rect 11885 16065 11897 16068
rect 11931 16096 11943 16099
rect 12406 16096 12434 16136
rect 15764 16108 15792 16136
rect 11931 16068 12434 16096
rect 11931 16065 11943 16068
rect 11885 16059 11943 16065
rect 15194 16056 15200 16108
rect 15252 16056 15258 16108
rect 15746 16056 15752 16108
rect 15804 16056 15810 16108
rect 21453 16099 21511 16105
rect 21453 16065 21465 16099
rect 21499 16065 21511 16099
rect 21560 16096 21588 16204
rect 21637 16201 21649 16235
rect 21683 16201 21695 16235
rect 21637 16195 21695 16201
rect 21652 16164 21680 16195
rect 21726 16192 21732 16244
rect 21784 16232 21790 16244
rect 23845 16235 23903 16241
rect 21784 16204 23520 16232
rect 21784 16192 21790 16204
rect 22066 16167 22124 16173
rect 22066 16164 22078 16167
rect 21652 16136 22078 16164
rect 22066 16133 22078 16136
rect 22112 16133 22124 16167
rect 23382 16164 23388 16176
rect 22066 16127 22124 16133
rect 23308 16136 23388 16164
rect 21560 16068 23152 16096
rect 21453 16059 21511 16065
rect 4798 15988 4804 16040
rect 4856 15988 4862 16040
rect 9692 16028 9720 16056
rect 10137 16031 10195 16037
rect 10137 16028 10149 16031
rect 9692 16000 10149 16028
rect 10137 15997 10149 16000
rect 10183 15997 10195 16031
rect 10137 15991 10195 15997
rect 10686 15988 10692 16040
rect 10744 16028 10750 16040
rect 10965 16031 11023 16037
rect 10965 16028 10977 16031
rect 10744 16000 10977 16028
rect 10744 15988 10750 16000
rect 10965 15997 10977 16000
rect 11011 15997 11023 16031
rect 10965 15991 11023 15997
rect 11057 16031 11115 16037
rect 11057 15997 11069 16031
rect 11103 15997 11115 16031
rect 15212 16028 15240 16056
rect 21358 16028 21364 16040
rect 15212 16000 21364 16028
rect 11057 15991 11115 15997
rect 9585 15963 9643 15969
rect 9585 15929 9597 15963
rect 9631 15960 9643 15963
rect 10045 15963 10103 15969
rect 10045 15960 10057 15963
rect 9631 15932 10057 15960
rect 9631 15929 9643 15932
rect 9585 15923 9643 15929
rect 10045 15929 10057 15932
rect 10091 15929 10103 15963
rect 10045 15923 10103 15929
rect 10413 15895 10471 15901
rect 10413 15861 10425 15895
rect 10459 15892 10471 15895
rect 10594 15892 10600 15904
rect 10459 15864 10600 15892
rect 10459 15861 10471 15864
rect 10413 15855 10471 15861
rect 10594 15852 10600 15864
rect 10652 15852 10658 15904
rect 10704 15892 10732 15988
rect 10778 15920 10784 15972
rect 10836 15960 10842 15972
rect 11072 15960 11100 15991
rect 21358 15988 21364 16000
rect 21416 15988 21422 16040
rect 10836 15932 11100 15960
rect 10836 15920 10842 15932
rect 15473 15895 15531 15901
rect 15473 15892 15485 15895
rect 10704 15864 15485 15892
rect 15473 15861 15485 15864
rect 15519 15892 15531 15895
rect 15562 15892 15568 15904
rect 15519 15864 15568 15892
rect 15519 15861 15531 15864
rect 15473 15855 15531 15861
rect 15562 15852 15568 15864
rect 15620 15852 15626 15904
rect 17954 15852 17960 15904
rect 18012 15892 18018 15904
rect 21174 15892 21180 15904
rect 18012 15864 21180 15892
rect 18012 15852 18018 15864
rect 21174 15852 21180 15864
rect 21232 15852 21238 15904
rect 21468 15892 21496 16059
rect 21542 15988 21548 16040
rect 21600 16028 21606 16040
rect 21821 16031 21879 16037
rect 21821 16028 21833 16031
rect 21600 16000 21833 16028
rect 21600 15988 21606 16000
rect 21821 15997 21833 16000
rect 21867 15997 21879 16031
rect 21821 15991 21879 15997
rect 22094 15892 22100 15904
rect 21468 15864 22100 15892
rect 22094 15852 22100 15864
rect 22152 15852 22158 15904
rect 23124 15892 23152 16068
rect 23198 16056 23204 16108
rect 23256 16056 23262 16108
rect 23308 16105 23336 16136
rect 23382 16124 23388 16136
rect 23440 16124 23446 16176
rect 23492 16173 23520 16204
rect 23845 16201 23857 16235
rect 23891 16232 23903 16235
rect 23891 16204 26004 16232
rect 23891 16201 23903 16204
rect 23845 16195 23903 16201
rect 23477 16167 23535 16173
rect 23477 16133 23489 16167
rect 23523 16133 23535 16167
rect 23477 16127 23535 16133
rect 23566 16124 23572 16176
rect 23624 16124 23630 16176
rect 25072 16167 25130 16173
rect 25072 16133 25084 16167
rect 25118 16164 25130 16167
rect 25866 16164 25872 16176
rect 25118 16136 25872 16164
rect 25118 16133 25130 16136
rect 25072 16127 25130 16133
rect 25866 16124 25872 16136
rect 25924 16124 25930 16176
rect 25976 16173 26004 16204
rect 26050 16192 26056 16244
rect 26108 16232 26114 16244
rect 27249 16235 27307 16241
rect 27249 16232 27261 16235
rect 26108 16204 27261 16232
rect 26108 16192 26114 16204
rect 27249 16201 27261 16204
rect 27295 16232 27307 16235
rect 27614 16232 27620 16244
rect 27295 16204 27620 16232
rect 27295 16201 27307 16204
rect 27249 16195 27307 16201
rect 27614 16192 27620 16204
rect 27672 16192 27678 16244
rect 25961 16167 26019 16173
rect 25961 16133 25973 16167
rect 26007 16133 26019 16167
rect 25961 16127 26019 16133
rect 23293 16099 23351 16105
rect 23293 16065 23305 16099
rect 23339 16065 23351 16099
rect 23293 16059 23351 16065
rect 23661 16099 23719 16105
rect 23661 16065 23673 16099
rect 23707 16065 23719 16099
rect 23661 16059 23719 16065
rect 25685 16099 25743 16105
rect 25685 16065 25697 16099
rect 25731 16065 25743 16099
rect 25685 16059 25743 16065
rect 23216 16028 23244 16056
rect 23676 16028 23704 16059
rect 23216 16000 23704 16028
rect 25317 16031 25375 16037
rect 25317 15997 25329 16031
rect 25363 16028 25375 16031
rect 25590 16028 25596 16040
rect 25363 16000 25596 16028
rect 25363 15997 25375 16000
rect 25317 15991 25375 15997
rect 25590 15988 25596 16000
rect 25648 15988 25654 16040
rect 25700 16028 25728 16059
rect 25774 16056 25780 16108
rect 25832 16056 25838 16108
rect 26142 16056 26148 16108
rect 26200 16096 26206 16108
rect 26329 16099 26387 16105
rect 26329 16096 26341 16099
rect 26200 16068 26341 16096
rect 26200 16056 26206 16068
rect 26329 16065 26341 16068
rect 26375 16065 26387 16099
rect 27154 16096 27160 16108
rect 26329 16059 26387 16065
rect 26436 16068 27160 16096
rect 26436 16028 26464 16068
rect 27154 16056 27160 16068
rect 27212 16056 27218 16108
rect 27341 16099 27399 16105
rect 27341 16065 27353 16099
rect 27387 16096 27399 16099
rect 27801 16099 27859 16105
rect 27801 16096 27813 16099
rect 27387 16068 27813 16096
rect 27387 16065 27399 16068
rect 27341 16059 27399 16065
rect 27801 16065 27813 16068
rect 27847 16065 27859 16099
rect 27801 16059 27859 16065
rect 25700 16000 26464 16028
rect 27062 15988 27068 16040
rect 27120 15988 27126 16040
rect 27890 15988 27896 16040
rect 27948 16028 27954 16040
rect 28353 16031 28411 16037
rect 28353 16028 28365 16031
rect 27948 16000 28365 16028
rect 27948 15988 27954 16000
rect 28353 15997 28365 16000
rect 28399 15997 28411 16031
rect 28353 15991 28411 15997
rect 23201 15963 23259 15969
rect 23201 15929 23213 15963
rect 23247 15960 23259 15963
rect 23566 15960 23572 15972
rect 23247 15932 23572 15960
rect 23247 15929 23259 15932
rect 23201 15923 23259 15929
rect 23566 15920 23572 15932
rect 23624 15920 23630 15972
rect 25501 15963 25559 15969
rect 23676 15932 24072 15960
rect 23676 15892 23704 15932
rect 23124 15864 23704 15892
rect 23934 15852 23940 15904
rect 23992 15852 23998 15904
rect 24044 15892 24072 15932
rect 25501 15929 25513 15963
rect 25547 15929 25559 15963
rect 25501 15923 25559 15929
rect 25516 15892 25544 15923
rect 24044 15864 25544 15892
rect 25961 15895 26019 15901
rect 25961 15861 25973 15895
rect 26007 15892 26019 15895
rect 26234 15892 26240 15904
rect 26007 15864 26240 15892
rect 26007 15861 26019 15864
rect 25961 15855 26019 15861
rect 26234 15852 26240 15864
rect 26292 15852 26298 15904
rect 26510 15852 26516 15904
rect 26568 15852 26574 15904
rect 27706 15852 27712 15904
rect 27764 15852 27770 15904
rect 1104 15802 31832 15824
rect 1104 15750 4182 15802
rect 4234 15750 4246 15802
rect 4298 15750 4310 15802
rect 4362 15750 4374 15802
rect 4426 15750 4438 15802
rect 4490 15750 4502 15802
rect 4554 15750 10182 15802
rect 10234 15750 10246 15802
rect 10298 15750 10310 15802
rect 10362 15750 10374 15802
rect 10426 15750 10438 15802
rect 10490 15750 10502 15802
rect 10554 15750 16182 15802
rect 16234 15750 16246 15802
rect 16298 15750 16310 15802
rect 16362 15750 16374 15802
rect 16426 15750 16438 15802
rect 16490 15750 16502 15802
rect 16554 15750 22182 15802
rect 22234 15750 22246 15802
rect 22298 15750 22310 15802
rect 22362 15750 22374 15802
rect 22426 15750 22438 15802
rect 22490 15750 22502 15802
rect 22554 15750 28182 15802
rect 28234 15750 28246 15802
rect 28298 15750 28310 15802
rect 28362 15750 28374 15802
rect 28426 15750 28438 15802
rect 28490 15750 28502 15802
rect 28554 15750 31832 15802
rect 1104 15728 31832 15750
rect 8297 15691 8355 15697
rect 8297 15657 8309 15691
rect 8343 15688 8355 15691
rect 8938 15688 8944 15700
rect 8343 15660 8944 15688
rect 8343 15657 8355 15660
rect 8297 15651 8355 15657
rect 8938 15648 8944 15660
rect 8996 15648 9002 15700
rect 9306 15648 9312 15700
rect 9364 15688 9370 15700
rect 10321 15691 10379 15697
rect 10321 15688 10333 15691
rect 9364 15660 10333 15688
rect 9364 15648 9370 15660
rect 10321 15657 10333 15660
rect 10367 15688 10379 15691
rect 10367 15660 11008 15688
rect 10367 15657 10379 15660
rect 10321 15651 10379 15657
rect 8754 15580 8760 15632
rect 8812 15580 8818 15632
rect 10980 15561 11008 15660
rect 15562 15648 15568 15700
rect 15620 15688 15626 15700
rect 22370 15688 22376 15700
rect 15620 15660 22376 15688
rect 15620 15648 15626 15660
rect 22370 15648 22376 15660
rect 22428 15648 22434 15700
rect 22465 15691 22523 15697
rect 22465 15657 22477 15691
rect 22511 15688 22523 15691
rect 22646 15688 22652 15700
rect 22511 15660 22652 15688
rect 22511 15657 22523 15660
rect 22465 15651 22523 15657
rect 22646 15648 22652 15660
rect 22704 15648 22710 15700
rect 23382 15648 23388 15700
rect 23440 15648 23446 15700
rect 26142 15648 26148 15700
rect 26200 15648 26206 15700
rect 27706 15648 27712 15700
rect 27764 15648 27770 15700
rect 21726 15620 21732 15632
rect 20640 15592 21732 15620
rect 8941 15555 8999 15561
rect 8941 15552 8953 15555
rect 8312 15524 8953 15552
rect 8312 15496 8340 15524
rect 8941 15521 8953 15524
rect 8987 15521 8999 15555
rect 8941 15515 8999 15521
rect 10965 15555 11023 15561
rect 10965 15521 10977 15555
rect 11011 15521 11023 15555
rect 10965 15515 11023 15521
rect 7190 15444 7196 15496
rect 7248 15484 7254 15496
rect 7745 15487 7803 15493
rect 7745 15484 7757 15487
rect 7248 15456 7757 15484
rect 7248 15444 7254 15456
rect 7745 15453 7757 15456
rect 7791 15453 7803 15487
rect 7745 15447 7803 15453
rect 7834 15444 7840 15496
rect 7892 15484 7898 15496
rect 8021 15487 8079 15493
rect 8021 15484 8033 15487
rect 7892 15456 8033 15484
rect 7892 15444 7898 15456
rect 8021 15453 8033 15456
rect 8067 15453 8079 15487
rect 8021 15447 8079 15453
rect 8113 15487 8171 15493
rect 8113 15453 8125 15487
rect 8159 15453 8171 15487
rect 8113 15447 8171 15453
rect 7929 15419 7987 15425
rect 7929 15385 7941 15419
rect 7975 15385 7987 15419
rect 8128 15416 8156 15447
rect 8294 15444 8300 15496
rect 8352 15444 8358 15496
rect 8570 15444 8576 15496
rect 8628 15444 8634 15496
rect 8680 15456 10272 15484
rect 8680 15416 8708 15456
rect 8128 15388 8708 15416
rect 7929 15379 7987 15385
rect 6638 15308 6644 15360
rect 6696 15308 6702 15360
rect 7944 15348 7972 15379
rect 8754 15376 8760 15428
rect 8812 15416 8818 15428
rect 9186 15419 9244 15425
rect 9186 15416 9198 15419
rect 8812 15388 9198 15416
rect 8812 15376 8818 15388
rect 9186 15385 9198 15388
rect 9232 15385 9244 15419
rect 10244 15416 10272 15456
rect 10410 15444 10416 15496
rect 10468 15444 10474 15496
rect 11974 15444 11980 15496
rect 12032 15444 12038 15496
rect 12621 15487 12679 15493
rect 12621 15453 12633 15487
rect 12667 15484 12679 15487
rect 12802 15484 12808 15496
rect 12667 15456 12808 15484
rect 12667 15453 12679 15456
rect 12621 15447 12679 15453
rect 12802 15444 12808 15456
rect 12860 15444 12866 15496
rect 17770 15444 17776 15496
rect 17828 15444 17834 15496
rect 18138 15444 18144 15496
rect 18196 15444 18202 15496
rect 18230 15444 18236 15496
rect 18288 15484 18294 15496
rect 18417 15487 18475 15493
rect 18417 15484 18429 15487
rect 18288 15456 18429 15484
rect 18288 15444 18294 15456
rect 18417 15453 18429 15456
rect 18463 15453 18475 15487
rect 18417 15447 18475 15453
rect 19889 15487 19947 15493
rect 19889 15453 19901 15487
rect 19935 15484 19947 15487
rect 20070 15484 20076 15496
rect 19935 15456 20076 15484
rect 19935 15453 19947 15456
rect 19889 15447 19947 15453
rect 20070 15444 20076 15456
rect 20128 15444 20134 15496
rect 20640 15493 20668 15592
rect 21726 15580 21732 15592
rect 21784 15580 21790 15632
rect 22554 15580 22560 15632
rect 22612 15620 22618 15632
rect 23198 15620 23204 15632
rect 22612 15592 23204 15620
rect 22612 15580 22618 15592
rect 23198 15580 23204 15592
rect 23256 15580 23262 15632
rect 20916 15524 21220 15552
rect 20916 15496 20944 15524
rect 20441 15487 20499 15493
rect 20441 15453 20453 15487
rect 20487 15453 20499 15487
rect 20441 15447 20499 15453
rect 20625 15487 20683 15493
rect 20625 15453 20637 15487
rect 20671 15453 20683 15487
rect 20625 15447 20683 15453
rect 20809 15487 20867 15493
rect 20809 15453 20821 15487
rect 20855 15484 20867 15487
rect 20898 15484 20904 15496
rect 20855 15456 20904 15484
rect 20855 15453 20867 15456
rect 20809 15447 20867 15453
rect 12526 15416 12532 15428
rect 10244 15388 12532 15416
rect 9186 15379 9244 15385
rect 12526 15376 12532 15388
rect 12584 15376 12590 15428
rect 18046 15376 18052 15428
rect 18104 15416 18110 15428
rect 19245 15419 19303 15425
rect 19245 15416 19257 15419
rect 18104 15388 19257 15416
rect 18104 15376 18110 15388
rect 19245 15385 19257 15388
rect 19291 15385 19303 15419
rect 19245 15379 19303 15385
rect 19702 15376 19708 15428
rect 19760 15416 19766 15428
rect 20456 15416 20484 15447
rect 20898 15444 20904 15456
rect 20956 15444 20962 15496
rect 20990 15444 20996 15496
rect 21048 15444 21054 15496
rect 21192 15484 21220 15524
rect 22922 15512 22928 15564
rect 22980 15512 22986 15564
rect 23014 15512 23020 15564
rect 23072 15512 23078 15564
rect 23400 15552 23428 15648
rect 23845 15555 23903 15561
rect 23845 15552 23857 15555
rect 23400 15524 23857 15552
rect 23845 15521 23857 15524
rect 23891 15521 23903 15555
rect 23845 15515 23903 15521
rect 25222 15512 25228 15564
rect 25280 15552 25286 15564
rect 25501 15555 25559 15561
rect 25501 15552 25513 15555
rect 25280 15524 25513 15552
rect 25280 15512 25286 15524
rect 25501 15521 25513 15524
rect 25547 15521 25559 15555
rect 27724 15552 27752 15648
rect 27724 15524 28672 15552
rect 25501 15515 25559 15521
rect 22462 15484 22468 15496
rect 21192 15456 22468 15484
rect 22462 15444 22468 15456
rect 22520 15444 22526 15496
rect 25590 15444 25596 15496
rect 25648 15484 25654 15496
rect 26237 15487 26295 15493
rect 26237 15484 26249 15487
rect 25648 15456 26249 15484
rect 25648 15444 25654 15456
rect 26237 15453 26249 15456
rect 26283 15484 26295 15487
rect 27522 15484 27528 15496
rect 26283 15456 27528 15484
rect 26283 15453 26295 15456
rect 26237 15447 26295 15453
rect 27522 15444 27528 15456
rect 27580 15444 27586 15496
rect 28644 15493 28672 15524
rect 28261 15487 28319 15493
rect 28261 15484 28273 15487
rect 27816 15456 28273 15484
rect 19760 15388 20484 15416
rect 20717 15419 20775 15425
rect 19760 15376 19766 15388
rect 20717 15385 20729 15419
rect 20763 15416 20775 15419
rect 21008 15416 21036 15444
rect 20763 15388 21036 15416
rect 22833 15419 22891 15425
rect 20763 15385 20775 15388
rect 20717 15379 20775 15385
rect 22833 15385 22845 15419
rect 22879 15416 22891 15419
rect 23293 15419 23351 15425
rect 23293 15416 23305 15419
rect 22879 15388 23305 15416
rect 22879 15385 22891 15388
rect 22833 15379 22891 15385
rect 23293 15385 23305 15388
rect 23339 15385 23351 15419
rect 23293 15379 23351 15385
rect 23934 15376 23940 15428
rect 23992 15416 23998 15428
rect 25685 15419 25743 15425
rect 25685 15416 25697 15419
rect 23992 15388 25697 15416
rect 23992 15376 23998 15388
rect 25685 15385 25697 15388
rect 25731 15416 25743 15419
rect 26050 15416 26056 15428
rect 25731 15388 26056 15416
rect 25731 15385 25743 15388
rect 25685 15379 25743 15385
rect 26050 15376 26056 15388
rect 26108 15376 26114 15428
rect 26510 15425 26516 15428
rect 26504 15416 26516 15425
rect 26471 15388 26516 15416
rect 26504 15379 26516 15388
rect 26510 15376 26516 15379
rect 26568 15376 26574 15428
rect 27709 15419 27767 15425
rect 27709 15416 27721 15419
rect 26712 15388 27721 15416
rect 12342 15348 12348 15360
rect 7944 15320 12348 15348
rect 12342 15308 12348 15320
rect 12400 15348 12406 15360
rect 12894 15348 12900 15360
rect 12400 15320 12900 15348
rect 12400 15308 12406 15320
rect 12894 15308 12900 15320
rect 12952 15308 12958 15360
rect 17586 15308 17592 15360
rect 17644 15308 17650 15360
rect 18325 15351 18383 15357
rect 18325 15317 18337 15351
rect 18371 15348 18383 15351
rect 18506 15348 18512 15360
rect 18371 15320 18512 15348
rect 18371 15317 18383 15320
rect 18325 15311 18383 15317
rect 18506 15308 18512 15320
rect 18564 15308 18570 15360
rect 18598 15308 18604 15360
rect 18656 15308 18662 15360
rect 20898 15308 20904 15360
rect 20956 15348 20962 15360
rect 20993 15351 21051 15357
rect 20993 15348 21005 15351
rect 20956 15320 21005 15348
rect 20956 15308 20962 15320
rect 20993 15317 21005 15320
rect 21039 15317 21051 15351
rect 20993 15311 21051 15317
rect 21174 15308 21180 15360
rect 21232 15348 21238 15360
rect 23014 15348 23020 15360
rect 21232 15320 23020 15348
rect 21232 15308 21238 15320
rect 23014 15308 23020 15320
rect 23072 15308 23078 15360
rect 25777 15351 25835 15357
rect 25777 15317 25789 15351
rect 25823 15348 25835 15351
rect 26712 15348 26740 15388
rect 27709 15385 27721 15388
rect 27755 15385 27767 15419
rect 27709 15379 27767 15385
rect 25823 15320 26740 15348
rect 25823 15317 25835 15320
rect 25777 15311 25835 15317
rect 27614 15308 27620 15360
rect 27672 15348 27678 15360
rect 27816 15348 27844 15456
rect 28261 15453 28273 15456
rect 28307 15453 28319 15487
rect 28261 15447 28319 15453
rect 28629 15487 28687 15493
rect 28629 15453 28641 15487
rect 28675 15453 28687 15487
rect 28629 15447 28687 15453
rect 27672 15320 27844 15348
rect 27672 15308 27678 15320
rect 28258 15308 28264 15360
rect 28316 15348 28322 15360
rect 28445 15351 28503 15357
rect 28445 15348 28457 15351
rect 28316 15320 28457 15348
rect 28316 15308 28322 15320
rect 28445 15317 28457 15320
rect 28491 15317 28503 15351
rect 28445 15311 28503 15317
rect 1104 15258 31832 15280
rect 1104 15206 4922 15258
rect 4974 15206 4986 15258
rect 5038 15206 5050 15258
rect 5102 15206 5114 15258
rect 5166 15206 5178 15258
rect 5230 15206 5242 15258
rect 5294 15206 10922 15258
rect 10974 15206 10986 15258
rect 11038 15206 11050 15258
rect 11102 15206 11114 15258
rect 11166 15206 11178 15258
rect 11230 15206 11242 15258
rect 11294 15206 16922 15258
rect 16974 15206 16986 15258
rect 17038 15206 17050 15258
rect 17102 15206 17114 15258
rect 17166 15206 17178 15258
rect 17230 15206 17242 15258
rect 17294 15206 22922 15258
rect 22974 15206 22986 15258
rect 23038 15206 23050 15258
rect 23102 15206 23114 15258
rect 23166 15206 23178 15258
rect 23230 15206 23242 15258
rect 23294 15206 28922 15258
rect 28974 15206 28986 15258
rect 29038 15206 29050 15258
rect 29102 15206 29114 15258
rect 29166 15206 29178 15258
rect 29230 15206 29242 15258
rect 29294 15206 31832 15258
rect 1104 15184 31832 15206
rect 3053 15147 3111 15153
rect 3053 15113 3065 15147
rect 3099 15113 3111 15147
rect 3053 15107 3111 15113
rect 2869 15011 2927 15017
rect 2869 14977 2881 15011
rect 2915 15008 2927 15011
rect 3068 15008 3096 15107
rect 6638 15104 6644 15156
rect 6696 15144 6702 15156
rect 6733 15147 6791 15153
rect 6733 15144 6745 15147
rect 6696 15116 6745 15144
rect 6696 15104 6702 15116
rect 6733 15113 6745 15116
rect 6779 15113 6791 15147
rect 6733 15107 6791 15113
rect 6822 15104 6828 15156
rect 6880 15104 6886 15156
rect 8021 15147 8079 15153
rect 8021 15113 8033 15147
rect 8067 15144 8079 15147
rect 8110 15144 8116 15156
rect 8067 15116 8116 15144
rect 8067 15113 8079 15116
rect 8021 15107 8079 15113
rect 8110 15104 8116 15116
rect 8168 15104 8174 15156
rect 8570 15104 8576 15156
rect 8628 15144 8634 15156
rect 8849 15147 8907 15153
rect 8849 15144 8861 15147
rect 8628 15116 8861 15144
rect 8628 15104 8634 15116
rect 8849 15113 8861 15116
rect 8895 15113 8907 15147
rect 8849 15107 8907 15113
rect 9217 15147 9275 15153
rect 9217 15113 9229 15147
rect 9263 15144 9275 15147
rect 10410 15144 10416 15156
rect 9263 15116 10416 15144
rect 9263 15113 9275 15116
rect 9217 15107 9275 15113
rect 10410 15104 10416 15116
rect 10468 15104 10474 15156
rect 12618 15104 12624 15156
rect 12676 15104 12682 15156
rect 18966 15104 18972 15156
rect 19024 15144 19030 15156
rect 19024 15116 21680 15144
rect 19024 15104 19030 15116
rect 8128 15076 8156 15104
rect 9309 15079 9367 15085
rect 9309 15076 9321 15079
rect 8128 15048 9321 15076
rect 9309 15045 9321 15048
rect 9355 15076 9367 15079
rect 10686 15076 10692 15088
rect 9355 15048 10692 15076
rect 9355 15045 9367 15048
rect 9309 15039 9367 15045
rect 10686 15036 10692 15048
rect 10744 15036 10750 15088
rect 12434 15085 12440 15088
rect 12428 15039 12440 15085
rect 12434 15036 12440 15039
rect 12492 15036 12498 15088
rect 12636 15076 12664 15104
rect 14642 15076 14648 15088
rect 12636 15048 14648 15076
rect 2915 14980 3096 15008
rect 3421 15011 3479 15017
rect 2915 14977 2927 14980
rect 2869 14971 2927 14977
rect 3421 14977 3433 15011
rect 3467 15008 3479 15011
rect 3881 15011 3939 15017
rect 3881 15008 3893 15011
rect 3467 14980 3893 15008
rect 3467 14977 3479 14980
rect 3421 14971 3479 14977
rect 3881 14977 3893 14980
rect 3927 14977 3939 15011
rect 3881 14971 3939 14977
rect 4448 14980 4844 15008
rect 1670 14900 1676 14952
rect 1728 14940 1734 14952
rect 3513 14943 3571 14949
rect 3513 14940 3525 14943
rect 1728 14912 3525 14940
rect 1728 14900 1734 14912
rect 3513 14909 3525 14912
rect 3559 14909 3571 14943
rect 3513 14903 3571 14909
rect 3697 14943 3755 14949
rect 3697 14909 3709 14943
rect 3743 14940 3755 14943
rect 4062 14940 4068 14952
rect 3743 14912 4068 14940
rect 3743 14909 3755 14912
rect 3697 14903 3755 14909
rect 3528 14816 3556 14903
rect 4062 14900 4068 14912
rect 4120 14940 4126 14952
rect 4448 14940 4476 14980
rect 4816 14952 4844 14980
rect 7926 14968 7932 15020
rect 7984 14968 7990 15020
rect 12636 15008 12664 15048
rect 14642 15036 14648 15048
rect 14700 15036 14706 15088
rect 18322 15076 18328 15088
rect 17328 15048 18328 15076
rect 9508 14980 12664 15008
rect 4120 14912 4476 14940
rect 4525 14943 4583 14949
rect 4120 14900 4126 14912
rect 4525 14909 4537 14943
rect 4571 14940 4583 14943
rect 4571 14912 4660 14940
rect 4571 14909 4583 14912
rect 4525 14903 4583 14909
rect 4632 14816 4660 14912
rect 4798 14900 4804 14952
rect 4856 14900 4862 14952
rect 7009 14943 7067 14949
rect 7009 14909 7021 14943
rect 7055 14940 7067 14943
rect 7098 14940 7104 14952
rect 7055 14912 7104 14940
rect 7055 14909 7067 14912
rect 7009 14903 7067 14909
rect 7098 14900 7104 14912
rect 7156 14900 7162 14952
rect 8202 14900 8208 14952
rect 8260 14900 8266 14952
rect 9508 14949 9536 14980
rect 13262 14968 13268 15020
rect 13320 15008 13326 15020
rect 17328 15017 17356 15048
rect 18322 15036 18328 15048
rect 18380 15076 18386 15088
rect 21542 15076 21548 15088
rect 18380 15048 21548 15076
rect 18380 15036 18386 15048
rect 17586 15017 17592 15020
rect 14921 15011 14979 15017
rect 14921 15008 14933 15011
rect 13320 14980 14933 15008
rect 13320 14968 13326 14980
rect 14921 14977 14933 14980
rect 14967 14977 14979 15011
rect 14921 14971 14979 14977
rect 17313 15011 17371 15017
rect 17313 14977 17325 15011
rect 17359 14977 17371 15011
rect 17580 15008 17592 15017
rect 17547 14980 17592 15008
rect 17313 14971 17371 14977
rect 17580 14971 17592 14980
rect 17586 14968 17592 14971
rect 17644 14968 17650 15020
rect 18506 14968 18512 15020
rect 18564 14968 18570 15020
rect 18800 15017 18828 15048
rect 21542 15036 21548 15048
rect 21600 15036 21606 15088
rect 21652 15076 21680 15116
rect 22094 15104 22100 15156
rect 22152 15144 22158 15156
rect 22189 15147 22247 15153
rect 22189 15144 22201 15147
rect 22152 15116 22201 15144
rect 22152 15104 22158 15116
rect 22189 15113 22201 15116
rect 22235 15113 22247 15147
rect 22189 15107 22247 15113
rect 22557 15147 22615 15153
rect 22557 15113 22569 15147
rect 22603 15144 22615 15147
rect 22738 15144 22744 15156
rect 22603 15116 22744 15144
rect 22603 15113 22615 15116
rect 22557 15107 22615 15113
rect 22738 15104 22744 15116
rect 22796 15104 22802 15156
rect 26234 15104 26240 15156
rect 26292 15104 26298 15156
rect 26973 15147 27031 15153
rect 26973 15113 26985 15147
rect 27019 15144 27031 15147
rect 27890 15144 27896 15156
rect 27019 15116 27896 15144
rect 27019 15113 27031 15116
rect 26973 15107 27031 15113
rect 26513 15079 26571 15085
rect 21652 15048 26372 15076
rect 18785 15011 18843 15017
rect 18785 14977 18797 15011
rect 18831 14977 18843 15011
rect 19041 15011 19099 15017
rect 19041 15008 19053 15011
rect 18785 14971 18843 14977
rect 18892 14980 19053 15008
rect 9493 14943 9551 14949
rect 9493 14909 9505 14943
rect 9539 14909 9551 14943
rect 9493 14903 9551 14909
rect 12161 14943 12219 14949
rect 12161 14909 12173 14943
rect 12207 14909 12219 14943
rect 14185 14943 14243 14949
rect 14185 14940 14197 14943
rect 12161 14903 12219 14909
rect 13556 14912 14197 14940
rect 2682 14764 2688 14816
rect 2740 14764 2746 14816
rect 3510 14764 3516 14816
rect 3568 14764 3574 14816
rect 4614 14764 4620 14816
rect 4672 14764 4678 14816
rect 6362 14764 6368 14816
rect 6420 14764 6426 14816
rect 7558 14764 7564 14816
rect 7616 14764 7622 14816
rect 12176 14804 12204 14903
rect 12526 14804 12532 14816
rect 12176 14776 12532 14804
rect 12526 14764 12532 14776
rect 12584 14764 12590 14816
rect 13446 14764 13452 14816
rect 13504 14804 13510 14816
rect 13556 14813 13584 14912
rect 14185 14909 14197 14912
rect 14231 14909 14243 14943
rect 18524 14940 18552 14968
rect 18892 14940 18920 14980
rect 19041 14977 19053 14980
rect 19087 14977 19099 15011
rect 19041 14971 19099 14977
rect 21266 14968 21272 15020
rect 21324 15008 21330 15020
rect 22005 15011 22063 15017
rect 22005 15008 22017 15011
rect 21324 14980 22017 15008
rect 21324 14968 21330 14980
rect 22005 14977 22017 14980
rect 22051 14977 22063 15011
rect 22005 14971 22063 14977
rect 22370 14968 22376 15020
rect 22428 15008 22434 15020
rect 22649 15011 22707 15017
rect 22649 15008 22661 15011
rect 22428 14980 22661 15008
rect 22428 14968 22434 14980
rect 22649 14977 22661 14980
rect 22695 15008 22707 15011
rect 23934 15008 23940 15020
rect 22695 14980 23940 15008
rect 22695 14977 22707 14980
rect 22649 14971 22707 14977
rect 23934 14968 23940 14980
rect 23992 14968 23998 15020
rect 20809 14943 20867 14949
rect 20809 14940 20821 14943
rect 18524 14912 18920 14940
rect 20180 14912 20821 14940
rect 14185 14903 14243 14909
rect 20180 14884 20208 14912
rect 20809 14909 20821 14912
rect 20855 14909 20867 14943
rect 20809 14903 20867 14909
rect 20990 14900 20996 14952
rect 21048 14900 21054 14952
rect 22741 14943 22799 14949
rect 21284 14912 22094 14940
rect 20162 14832 20168 14884
rect 20220 14832 20226 14884
rect 21284 14872 21312 14912
rect 20824 14844 21312 14872
rect 20824 14816 20852 14844
rect 21358 14832 21364 14884
rect 21416 14872 21422 14884
rect 21821 14875 21879 14881
rect 21821 14872 21833 14875
rect 21416 14844 21833 14872
rect 21416 14832 21422 14844
rect 21821 14841 21833 14844
rect 21867 14841 21879 14875
rect 22066 14872 22094 14912
rect 22741 14909 22753 14943
rect 22787 14909 22799 14943
rect 22741 14903 22799 14909
rect 22756 14872 22784 14903
rect 22066 14844 22784 14872
rect 21821 14835 21879 14841
rect 13541 14807 13599 14813
rect 13541 14804 13553 14807
rect 13504 14776 13553 14804
rect 13504 14764 13510 14776
rect 13541 14773 13553 14776
rect 13587 14773 13599 14807
rect 13541 14767 13599 14773
rect 13630 14764 13636 14816
rect 13688 14764 13694 14816
rect 14366 14764 14372 14816
rect 14424 14764 14430 14816
rect 18693 14807 18751 14813
rect 18693 14773 18705 14807
rect 18739 14804 18751 14807
rect 20070 14804 20076 14816
rect 18739 14776 20076 14804
rect 18739 14773 18751 14776
rect 18693 14767 18751 14773
rect 20070 14764 20076 14776
rect 20128 14764 20134 14816
rect 20254 14764 20260 14816
rect 20312 14764 20318 14816
rect 20806 14764 20812 14816
rect 20864 14764 20870 14816
rect 21634 14764 21640 14816
rect 21692 14764 21698 14816
rect 26344 14804 26372 15048
rect 26513 15045 26525 15079
rect 26559 15076 26571 15079
rect 26988 15076 27016 15107
rect 27890 15104 27896 15116
rect 27948 15104 27954 15156
rect 26559 15048 27016 15076
rect 26559 15045 26571 15048
rect 26513 15039 26571 15045
rect 27522 15036 27528 15088
rect 27580 15076 27586 15088
rect 27580 15048 28396 15076
rect 27580 15036 27586 15048
rect 26418 14968 26424 15020
rect 26476 14968 26482 15020
rect 26605 15011 26663 15017
rect 26605 14977 26617 15011
rect 26651 15008 26663 15011
rect 26694 15008 26700 15020
rect 26651 14980 26700 15008
rect 26651 14977 26663 14980
rect 26605 14971 26663 14977
rect 26694 14968 26700 14980
rect 26752 14968 26758 15020
rect 26789 15011 26847 15017
rect 26789 14977 26801 15011
rect 26835 15008 26847 15011
rect 27614 15008 27620 15020
rect 26835 14980 27620 15008
rect 26835 14977 26847 14980
rect 26789 14971 26847 14977
rect 27614 14968 27620 14980
rect 27672 14968 27678 15020
rect 28097 15011 28155 15017
rect 28097 14977 28109 15011
rect 28143 15008 28155 15011
rect 28258 15008 28264 15020
rect 28143 14980 28264 15008
rect 28143 14977 28155 14980
rect 28097 14971 28155 14977
rect 28258 14968 28264 14980
rect 28316 14968 28322 15020
rect 28368 15017 28396 15048
rect 28353 15011 28411 15017
rect 28353 14977 28365 15011
rect 28399 15008 28411 15011
rect 28626 15008 28632 15020
rect 28399 14980 28632 15008
rect 28399 14977 28411 14980
rect 28353 14971 28411 14977
rect 28626 14968 28632 14980
rect 28684 14968 28690 15020
rect 31202 14804 31208 14816
rect 26344 14776 31208 14804
rect 31202 14764 31208 14776
rect 31260 14764 31266 14816
rect 1104 14714 31832 14736
rect 1104 14662 4182 14714
rect 4234 14662 4246 14714
rect 4298 14662 4310 14714
rect 4362 14662 4374 14714
rect 4426 14662 4438 14714
rect 4490 14662 4502 14714
rect 4554 14662 10182 14714
rect 10234 14662 10246 14714
rect 10298 14662 10310 14714
rect 10362 14662 10374 14714
rect 10426 14662 10438 14714
rect 10490 14662 10502 14714
rect 10554 14662 16182 14714
rect 16234 14662 16246 14714
rect 16298 14662 16310 14714
rect 16362 14662 16374 14714
rect 16426 14662 16438 14714
rect 16490 14662 16502 14714
rect 16554 14662 22182 14714
rect 22234 14662 22246 14714
rect 22298 14662 22310 14714
rect 22362 14662 22374 14714
rect 22426 14662 22438 14714
rect 22490 14662 22502 14714
rect 22554 14662 28182 14714
rect 28234 14662 28246 14714
rect 28298 14662 28310 14714
rect 28362 14662 28374 14714
rect 28426 14662 28438 14714
rect 28490 14662 28502 14714
rect 28554 14662 31832 14714
rect 1104 14640 31832 14662
rect 6365 14603 6423 14609
rect 6365 14569 6377 14603
rect 6411 14600 6423 14603
rect 7190 14600 7196 14612
rect 6411 14572 7196 14600
rect 6411 14569 6423 14572
rect 6365 14563 6423 14569
rect 7190 14560 7196 14572
rect 7248 14560 7254 14612
rect 7834 14560 7840 14612
rect 7892 14560 7898 14612
rect 7926 14560 7932 14612
rect 7984 14560 7990 14612
rect 12434 14560 12440 14612
rect 12492 14560 12498 14612
rect 13630 14560 13636 14612
rect 13688 14560 13694 14612
rect 17770 14560 17776 14612
rect 17828 14600 17834 14612
rect 17865 14603 17923 14609
rect 17865 14600 17877 14603
rect 17828 14572 17877 14600
rect 17828 14560 17834 14572
rect 17865 14569 17877 14572
rect 17911 14569 17923 14603
rect 17865 14563 17923 14569
rect 17954 14560 17960 14612
rect 18012 14560 18018 14612
rect 18138 14560 18144 14612
rect 18196 14600 18202 14612
rect 19245 14603 19303 14609
rect 19245 14600 19257 14603
rect 18196 14572 19257 14600
rect 18196 14560 18202 14572
rect 19245 14569 19257 14572
rect 19291 14569 19303 14603
rect 20254 14600 20260 14612
rect 19245 14563 19303 14569
rect 19628 14572 20260 14600
rect 12713 14535 12771 14541
rect 12713 14501 12725 14535
rect 12759 14501 12771 14535
rect 12713 14495 12771 14501
rect 4433 14467 4491 14473
rect 4433 14433 4445 14467
rect 4479 14464 4491 14467
rect 4706 14464 4712 14476
rect 4479 14436 4712 14464
rect 4479 14433 4491 14436
rect 4433 14427 4491 14433
rect 4706 14424 4712 14436
rect 4764 14424 4770 14476
rect 10597 14467 10655 14473
rect 10597 14464 10609 14467
rect 8312 14436 10609 14464
rect 8312 14408 8340 14436
rect 10597 14433 10609 14436
rect 10643 14433 10655 14467
rect 10597 14427 10655 14433
rect 2225 14399 2283 14405
rect 2225 14365 2237 14399
rect 2271 14396 2283 14399
rect 4985 14399 5043 14405
rect 4985 14396 4997 14399
rect 2271 14368 4997 14396
rect 2271 14365 2283 14368
rect 2225 14359 2283 14365
rect 2332 14272 2360 14368
rect 4985 14365 4997 14368
rect 5031 14396 5043 14399
rect 6457 14399 6515 14405
rect 6457 14396 6469 14399
rect 5031 14368 6469 14396
rect 5031 14365 5043 14368
rect 4985 14359 5043 14365
rect 6457 14365 6469 14368
rect 6503 14396 6515 14399
rect 8294 14396 8300 14408
rect 6503 14368 8300 14396
rect 6503 14365 6515 14368
rect 6457 14359 6515 14365
rect 8294 14356 8300 14368
rect 8352 14356 8358 14408
rect 8481 14399 8539 14405
rect 8481 14365 8493 14399
rect 8527 14365 8539 14399
rect 12621 14399 12679 14405
rect 8481 14359 8539 14365
rect 8588 14368 11928 14396
rect 2492 14331 2550 14337
rect 2492 14297 2504 14331
rect 2538 14328 2550 14331
rect 3234 14328 3240 14340
rect 2538 14300 3240 14328
rect 2538 14297 2550 14300
rect 2492 14291 2550 14297
rect 3234 14288 3240 14300
rect 3292 14288 3298 14340
rect 3510 14288 3516 14340
rect 3568 14328 3574 14340
rect 5252 14331 5310 14337
rect 3568 14300 4292 14328
rect 3568 14288 3574 14300
rect 2314 14220 2320 14272
rect 2372 14220 2378 14272
rect 3602 14220 3608 14272
rect 3660 14220 3666 14272
rect 3786 14220 3792 14272
rect 3844 14220 3850 14272
rect 4154 14220 4160 14272
rect 4212 14220 4218 14272
rect 4264 14269 4292 14300
rect 5252 14297 5264 14331
rect 5298 14328 5310 14331
rect 5994 14328 6000 14340
rect 5298 14300 6000 14328
rect 5298 14297 5310 14300
rect 5252 14291 5310 14297
rect 5994 14288 6000 14300
rect 6052 14288 6058 14340
rect 6724 14331 6782 14337
rect 6724 14297 6736 14331
rect 6770 14328 6782 14331
rect 7006 14328 7012 14340
rect 6770 14300 7012 14328
rect 6770 14297 6782 14300
rect 6724 14291 6782 14297
rect 7006 14288 7012 14300
rect 7064 14288 7070 14340
rect 7834 14288 7840 14340
rect 7892 14328 7898 14340
rect 8496 14328 8524 14359
rect 7892 14300 8524 14328
rect 7892 14288 7898 14300
rect 4249 14263 4307 14269
rect 4249 14229 4261 14263
rect 4295 14260 4307 14263
rect 8588 14260 8616 14368
rect 10864 14331 10922 14337
rect 10864 14297 10876 14331
rect 10910 14297 10922 14331
rect 10864 14291 10922 14297
rect 11900 14328 11928 14368
rect 12621 14365 12633 14399
rect 12667 14396 12679 14399
rect 12728 14396 12756 14495
rect 13354 14424 13360 14476
rect 13412 14464 13418 14476
rect 13538 14464 13544 14476
rect 13412 14436 13544 14464
rect 13412 14424 13418 14436
rect 13538 14424 13544 14436
rect 13596 14424 13602 14476
rect 12667 14368 12756 14396
rect 13081 14399 13139 14405
rect 12667 14365 12679 14368
rect 12621 14359 12679 14365
rect 13081 14365 13093 14399
rect 13127 14396 13139 14399
rect 13648 14396 13676 14560
rect 16022 14492 16028 14544
rect 16080 14532 16086 14544
rect 17972 14532 18000 14560
rect 16080 14504 16712 14532
rect 16080 14492 16086 14504
rect 16684 14473 16712 14504
rect 17236 14504 18000 14532
rect 17236 14473 17264 14504
rect 14645 14467 14703 14473
rect 14645 14464 14657 14467
rect 14108 14436 14657 14464
rect 14108 14408 14136 14436
rect 14645 14433 14657 14436
rect 14691 14433 14703 14467
rect 14645 14427 14703 14433
rect 16669 14467 16727 14473
rect 16669 14433 16681 14467
rect 16715 14433 16727 14467
rect 16669 14427 16727 14433
rect 17221 14467 17279 14473
rect 17221 14433 17233 14467
rect 17267 14433 17279 14467
rect 18325 14467 18383 14473
rect 18325 14464 18337 14467
rect 17221 14427 17279 14433
rect 17328 14436 18337 14464
rect 13127 14368 13676 14396
rect 13127 14365 13139 14368
rect 13081 14359 13139 14365
rect 13722 14356 13728 14408
rect 13780 14356 13786 14408
rect 14090 14356 14096 14408
rect 14148 14356 14154 14408
rect 14369 14399 14427 14405
rect 14369 14365 14381 14399
rect 14415 14396 14427 14399
rect 14734 14396 14740 14408
rect 14415 14368 14740 14396
rect 14415 14365 14427 14368
rect 14369 14359 14427 14365
rect 14734 14356 14740 14368
rect 14792 14356 14798 14408
rect 13173 14331 13231 14337
rect 13173 14328 13185 14331
rect 11900 14300 13185 14328
rect 4295 14232 8616 14260
rect 4295 14229 4307 14232
rect 4249 14223 4307 14229
rect 10778 14220 10784 14272
rect 10836 14260 10842 14272
rect 10888 14260 10916 14291
rect 11900 14272 11928 14300
rect 13173 14297 13185 14300
rect 13219 14328 13231 14331
rect 14458 14328 14464 14340
rect 13219 14300 14464 14328
rect 13219 14297 13231 14300
rect 13173 14291 13231 14297
rect 14458 14288 14464 14300
rect 14516 14288 14522 14340
rect 14890 14331 14948 14337
rect 14890 14328 14902 14331
rect 14568 14300 14902 14328
rect 10836 14232 10916 14260
rect 10836 14220 10842 14232
rect 11882 14220 11888 14272
rect 11940 14220 11946 14272
rect 11977 14263 12035 14269
rect 11977 14229 11989 14263
rect 12023 14260 12035 14263
rect 12802 14260 12808 14272
rect 12023 14232 12808 14260
rect 12023 14229 12035 14232
rect 11977 14223 12035 14229
rect 12802 14220 12808 14232
rect 12860 14220 12866 14272
rect 13538 14220 13544 14272
rect 13596 14220 13602 14272
rect 14568 14269 14596 14300
rect 14890 14297 14902 14300
rect 14936 14297 14948 14331
rect 14890 14291 14948 14297
rect 14553 14263 14611 14269
rect 14553 14229 14565 14263
rect 14599 14229 14611 14263
rect 14553 14223 14611 14229
rect 16114 14220 16120 14272
rect 16172 14220 16178 14272
rect 16666 14220 16672 14272
rect 16724 14260 16730 14272
rect 17328 14269 17356 14436
rect 18325 14433 18337 14436
rect 18371 14433 18383 14467
rect 18325 14427 18383 14433
rect 18506 14424 18512 14476
rect 18564 14464 18570 14476
rect 19150 14464 19156 14476
rect 18564 14436 19156 14464
rect 18564 14424 18570 14436
rect 19150 14424 19156 14436
rect 19208 14424 19214 14476
rect 17405 14399 17463 14405
rect 17405 14365 17417 14399
rect 17451 14396 17463 14399
rect 18138 14396 18144 14408
rect 17451 14368 18144 14396
rect 17451 14365 17463 14368
rect 17405 14359 17463 14365
rect 18138 14356 18144 14368
rect 18196 14356 18202 14408
rect 18230 14356 18236 14408
rect 18288 14356 18294 14408
rect 19628 14405 19656 14572
rect 20254 14560 20260 14572
rect 20312 14560 20318 14612
rect 20898 14560 20904 14612
rect 20956 14600 20962 14612
rect 21726 14600 21732 14612
rect 20956 14572 21732 14600
rect 20956 14560 20962 14572
rect 21726 14560 21732 14572
rect 21784 14560 21790 14612
rect 19886 14424 19892 14476
rect 19944 14424 19950 14476
rect 19613 14399 19671 14405
rect 19613 14365 19625 14399
rect 19659 14365 19671 14399
rect 19613 14359 19671 14365
rect 21358 14356 21364 14408
rect 21416 14405 21422 14408
rect 21416 14396 21428 14405
rect 21416 14368 21461 14396
rect 21416 14359 21428 14368
rect 21416 14356 21422 14359
rect 21542 14356 21548 14408
rect 21600 14396 21606 14408
rect 21637 14399 21695 14405
rect 21637 14396 21649 14399
rect 21600 14368 21649 14396
rect 21600 14356 21606 14368
rect 21637 14365 21649 14368
rect 21683 14365 21695 14399
rect 21637 14359 21695 14365
rect 18248 14328 18276 14356
rect 17788 14300 18276 14328
rect 19705 14331 19763 14337
rect 17788 14269 17816 14300
rect 19705 14297 19717 14331
rect 19751 14328 19763 14331
rect 19751 14300 21128 14328
rect 19751 14297 19763 14300
rect 19705 14291 19763 14297
rect 21100 14272 21128 14300
rect 17313 14263 17371 14269
rect 17313 14260 17325 14263
rect 16724 14232 17325 14260
rect 16724 14220 16730 14232
rect 17313 14229 17325 14232
rect 17359 14229 17371 14263
rect 17313 14223 17371 14229
rect 17773 14263 17831 14269
rect 17773 14229 17785 14263
rect 17819 14229 17831 14263
rect 17773 14223 17831 14229
rect 18046 14220 18052 14272
rect 18104 14260 18110 14272
rect 18233 14263 18291 14269
rect 18233 14260 18245 14263
rect 18104 14232 18245 14260
rect 18104 14220 18110 14232
rect 18233 14229 18245 14232
rect 18279 14229 18291 14263
rect 18233 14223 18291 14229
rect 20257 14263 20315 14269
rect 20257 14229 20269 14263
rect 20303 14260 20315 14263
rect 20990 14260 20996 14272
rect 20303 14232 20996 14260
rect 20303 14229 20315 14232
rect 20257 14223 20315 14229
rect 20990 14220 20996 14232
rect 21048 14220 21054 14272
rect 21082 14220 21088 14272
rect 21140 14220 21146 14272
rect 1104 14170 31832 14192
rect 1104 14118 4922 14170
rect 4974 14118 4986 14170
rect 5038 14118 5050 14170
rect 5102 14118 5114 14170
rect 5166 14118 5178 14170
rect 5230 14118 5242 14170
rect 5294 14118 10922 14170
rect 10974 14118 10986 14170
rect 11038 14118 11050 14170
rect 11102 14118 11114 14170
rect 11166 14118 11178 14170
rect 11230 14118 11242 14170
rect 11294 14118 16922 14170
rect 16974 14118 16986 14170
rect 17038 14118 17050 14170
rect 17102 14118 17114 14170
rect 17166 14118 17178 14170
rect 17230 14118 17242 14170
rect 17294 14118 22922 14170
rect 22974 14118 22986 14170
rect 23038 14118 23050 14170
rect 23102 14118 23114 14170
rect 23166 14118 23178 14170
rect 23230 14118 23242 14170
rect 23294 14118 28922 14170
rect 28974 14118 28986 14170
rect 29038 14118 29050 14170
rect 29102 14118 29114 14170
rect 29166 14118 29178 14170
rect 29230 14118 29242 14170
rect 29294 14118 31832 14170
rect 1104 14096 31832 14118
rect 2682 14016 2688 14068
rect 2740 14016 2746 14068
rect 3602 14016 3608 14068
rect 3660 14016 3666 14068
rect 3697 14059 3755 14065
rect 3697 14025 3709 14059
rect 3743 14025 3755 14059
rect 3697 14019 3755 14025
rect 3973 14059 4031 14065
rect 3973 14025 3985 14059
rect 4019 14056 4031 14059
rect 4154 14056 4160 14068
rect 4019 14028 4160 14056
rect 4019 14025 4031 14028
rect 3973 14019 4031 14025
rect 2584 13991 2642 13997
rect 2584 13957 2596 13991
rect 2630 13988 2642 13991
rect 2700 13988 2728 14016
rect 2630 13960 2728 13988
rect 2630 13957 2642 13960
rect 2584 13951 2642 13957
rect 2314 13880 2320 13932
rect 2372 13880 2378 13932
rect 3620 13920 3648 14016
rect 3712 13988 3740 14019
rect 4154 14016 4160 14028
rect 4212 14016 4218 14068
rect 5350 14056 5356 14068
rect 5092 14028 5356 14056
rect 4614 13988 4620 14000
rect 3712 13960 4620 13988
rect 4614 13948 4620 13960
rect 4672 13988 4678 14000
rect 4985 13991 5043 13997
rect 4985 13988 4997 13991
rect 4672 13960 4997 13988
rect 4672 13948 4678 13960
rect 4985 13957 4997 13960
rect 5031 13957 5043 13991
rect 4985 13951 5043 13957
rect 5092 13929 5120 14028
rect 5350 14016 5356 14028
rect 5408 14056 5414 14068
rect 5810 14056 5816 14068
rect 5408 14028 5816 14056
rect 5408 14016 5414 14028
rect 5810 14016 5816 14028
rect 5868 14016 5874 14068
rect 5994 14016 6000 14068
rect 6052 14016 6058 14068
rect 6362 14016 6368 14068
rect 6420 14016 6426 14068
rect 7006 14016 7012 14068
rect 7064 14016 7070 14068
rect 7558 14016 7564 14068
rect 7616 14016 7622 14068
rect 10778 14016 10784 14068
rect 10836 14056 10842 14068
rect 10965 14059 11023 14065
rect 10965 14056 10977 14059
rect 10836 14028 10977 14056
rect 10836 14016 10842 14028
rect 10965 14025 10977 14028
rect 11011 14025 11023 14059
rect 10965 14019 11023 14025
rect 11517 14059 11575 14065
rect 11517 14025 11529 14059
rect 11563 14025 11575 14059
rect 11517 14019 11575 14025
rect 11885 14059 11943 14065
rect 11885 14025 11897 14059
rect 11931 14056 11943 14059
rect 11974 14056 11980 14068
rect 11931 14028 11980 14056
rect 11931 14025 11943 14028
rect 11885 14019 11943 14025
rect 5442 13988 5448 14000
rect 5184 13960 5448 13988
rect 4525 13923 4583 13929
rect 4525 13920 4537 13923
rect 3620 13892 4537 13920
rect 4525 13889 4537 13892
rect 4571 13920 4583 13923
rect 4709 13923 4767 13929
rect 4709 13920 4721 13923
rect 4571 13892 4721 13920
rect 4571 13889 4583 13892
rect 4525 13883 4583 13889
rect 4709 13889 4721 13892
rect 4755 13889 4767 13923
rect 4709 13883 4767 13889
rect 4893 13923 4951 13929
rect 4893 13889 4905 13923
rect 4939 13889 4951 13923
rect 4893 13883 4951 13889
rect 5077 13923 5135 13929
rect 5077 13889 5089 13923
rect 5123 13889 5135 13923
rect 5077 13883 5135 13889
rect 4908 13852 4936 13883
rect 5184 13852 5212 13960
rect 5442 13948 5448 13960
rect 5500 13988 5506 14000
rect 5718 13988 5724 14000
rect 5500 13960 5724 13988
rect 5500 13948 5506 13960
rect 5718 13948 5724 13960
rect 5776 13948 5782 14000
rect 6181 13923 6239 13929
rect 6181 13889 6193 13923
rect 6227 13920 6239 13923
rect 6380 13920 6408 14016
rect 6227 13892 6408 13920
rect 7193 13923 7251 13929
rect 6227 13889 6239 13892
rect 6181 13883 6239 13889
rect 7193 13889 7205 13923
rect 7239 13920 7251 13923
rect 7576 13920 7604 14016
rect 7239 13892 7604 13920
rect 11149 13923 11207 13929
rect 7239 13889 7251 13892
rect 7193 13883 7251 13889
rect 11149 13889 11161 13923
rect 11195 13920 11207 13923
rect 11532 13920 11560 14019
rect 11974 14016 11980 14028
rect 12032 14016 12038 14068
rect 12437 14059 12495 14065
rect 12437 14025 12449 14059
rect 12483 14056 12495 14059
rect 13078 14056 13084 14068
rect 12483 14028 13084 14056
rect 12483 14025 12495 14028
rect 12437 14019 12495 14025
rect 13078 14016 13084 14028
rect 13136 14056 13142 14068
rect 13262 14056 13268 14068
rect 13136 14028 13268 14056
rect 13136 14016 13142 14028
rect 13262 14016 13268 14028
rect 13320 14016 13326 14068
rect 13722 14016 13728 14068
rect 13780 14056 13786 14068
rect 13909 14059 13967 14065
rect 13909 14056 13921 14059
rect 13780 14028 13921 14056
rect 13780 14016 13786 14028
rect 13909 14025 13921 14028
rect 13955 14025 13967 14059
rect 13909 14019 13967 14025
rect 14277 14059 14335 14065
rect 14277 14025 14289 14059
rect 14323 14056 14335 14059
rect 14366 14056 14372 14068
rect 14323 14028 14372 14056
rect 14323 14025 14335 14028
rect 14277 14019 14335 14025
rect 14366 14016 14372 14028
rect 14424 14016 14430 14068
rect 14458 14016 14464 14068
rect 14516 14016 14522 14068
rect 14734 14016 14740 14068
rect 14792 14056 14798 14068
rect 14921 14059 14979 14065
rect 14921 14056 14933 14059
rect 14792 14028 14933 14056
rect 14792 14016 14798 14028
rect 14921 14025 14933 14028
rect 14967 14025 14979 14059
rect 14921 14019 14979 14025
rect 15289 14059 15347 14065
rect 15289 14025 15301 14059
rect 15335 14056 15347 14059
rect 16114 14056 16120 14068
rect 15335 14028 16120 14056
rect 15335 14025 15347 14028
rect 15289 14019 15347 14025
rect 16114 14016 16120 14028
rect 16172 14016 16178 14068
rect 18322 14016 18328 14068
rect 18380 14016 18386 14068
rect 19702 14016 19708 14068
rect 19760 14016 19766 14068
rect 20162 14056 20168 14068
rect 19812 14028 20168 14056
rect 13538 13948 13544 14000
rect 13596 13997 13602 14000
rect 13596 13988 13608 13997
rect 14476 13988 14504 14016
rect 15933 13991 15991 13997
rect 13596 13960 13641 13988
rect 14476 13960 15884 13988
rect 13596 13951 13608 13960
rect 13596 13948 13602 13951
rect 11195 13892 11560 13920
rect 11624 13892 15700 13920
rect 11195 13889 11207 13892
rect 11149 13883 11207 13889
rect 11624 13852 11652 13892
rect 4908 13824 5212 13852
rect 5276 13824 11652 13852
rect 5276 13793 5304 13824
rect 11882 13812 11888 13864
rect 11940 13852 11946 13864
rect 11977 13855 12035 13861
rect 11977 13852 11989 13855
rect 11940 13824 11989 13852
rect 11940 13812 11946 13824
rect 11977 13821 11989 13824
rect 12023 13821 12035 13855
rect 11977 13815 12035 13821
rect 12066 13812 12072 13864
rect 12124 13812 12130 13864
rect 13817 13855 13875 13861
rect 13817 13821 13829 13855
rect 13863 13852 13875 13855
rect 14090 13852 14096 13864
rect 13863 13824 14096 13852
rect 13863 13821 13875 13824
rect 13817 13815 13875 13821
rect 14090 13812 14096 13824
rect 14148 13812 14154 13864
rect 14369 13855 14427 13861
rect 14369 13821 14381 13855
rect 14415 13821 14427 13855
rect 14369 13815 14427 13821
rect 5261 13787 5319 13793
rect 5261 13753 5273 13787
rect 5307 13753 5319 13787
rect 14384 13784 14412 13815
rect 14458 13812 14464 13864
rect 14516 13812 14522 13864
rect 15378 13852 15384 13864
rect 14568 13824 15384 13852
rect 14568 13796 14596 13824
rect 15378 13812 15384 13824
rect 15436 13812 15442 13864
rect 15565 13855 15623 13861
rect 15565 13821 15577 13855
rect 15611 13821 15623 13855
rect 15672 13852 15700 13892
rect 15746 13880 15752 13932
rect 15804 13880 15810 13932
rect 15856 13920 15884 13960
rect 15933 13957 15945 13991
rect 15979 13988 15991 13991
rect 16022 13988 16028 14000
rect 15979 13960 16028 13988
rect 15979 13957 15991 13960
rect 15933 13951 15991 13957
rect 16022 13948 16028 13960
rect 16080 13948 16086 14000
rect 16666 13920 16672 13932
rect 15856 13892 16672 13920
rect 16666 13880 16672 13892
rect 16724 13880 16730 13932
rect 18340 13929 18368 14016
rect 18598 13997 18604 14000
rect 18592 13988 18604 13997
rect 18559 13960 18604 13988
rect 18592 13951 18604 13960
rect 18598 13948 18604 13951
rect 18656 13948 18662 14000
rect 19812 13929 19840 14028
rect 20162 14016 20168 14028
rect 20220 14016 20226 14068
rect 20254 14016 20260 14068
rect 20312 14016 20318 14068
rect 20349 14059 20407 14065
rect 20349 14025 20361 14059
rect 20395 14025 20407 14059
rect 20349 14019 20407 14025
rect 21085 14059 21143 14065
rect 21085 14025 21097 14059
rect 21131 14056 21143 14059
rect 21634 14056 21640 14068
rect 21131 14028 21640 14056
rect 21131 14025 21143 14028
rect 21085 14019 21143 14025
rect 19978 13948 19984 14000
rect 20036 13948 20042 14000
rect 20070 13948 20076 14000
rect 20128 13948 20134 14000
rect 20272 13988 20300 14016
rect 20180 13960 20300 13988
rect 20364 13988 20392 14019
rect 21634 14016 21640 14028
rect 21692 14016 21698 14068
rect 22094 14016 22100 14068
rect 22152 14056 22158 14068
rect 22281 14059 22339 14065
rect 22281 14056 22293 14059
rect 22152 14028 22293 14056
rect 22152 14016 22158 14028
rect 22281 14025 22293 14028
rect 22327 14025 22339 14059
rect 26418 14056 26424 14068
rect 22281 14019 22339 14025
rect 24964 14028 26424 14056
rect 20364 13960 22048 13988
rect 20180 13929 20208 13960
rect 18325 13923 18383 13929
rect 18325 13889 18337 13923
rect 18371 13889 18383 13923
rect 19797 13923 19855 13929
rect 18325 13883 18383 13889
rect 18432 13892 19380 13920
rect 16574 13852 16580 13864
rect 15672 13824 16580 13852
rect 15565 13815 15623 13821
rect 14550 13784 14556 13796
rect 14384 13756 14556 13784
rect 5261 13747 5319 13753
rect 14550 13744 14556 13756
rect 14608 13744 14614 13796
rect 14918 13744 14924 13796
rect 14976 13784 14982 13796
rect 15580 13784 15608 13815
rect 16574 13812 16580 13824
rect 16632 13812 16638 13864
rect 18432 13852 18460 13892
rect 16868 13824 18460 13852
rect 19352 13852 19380 13892
rect 19797 13889 19809 13923
rect 19843 13889 19855 13923
rect 19797 13883 19855 13889
rect 20165 13923 20223 13929
rect 20165 13889 20177 13923
rect 20211 13889 20223 13923
rect 20993 13923 21051 13929
rect 20993 13920 21005 13923
rect 20165 13883 20223 13889
rect 20272 13892 21005 13920
rect 20272 13852 20300 13892
rect 20993 13889 21005 13892
rect 21039 13920 21051 13923
rect 21082 13920 21088 13932
rect 21039 13892 21088 13920
rect 21039 13889 21051 13892
rect 20993 13883 21051 13889
rect 21082 13880 21088 13892
rect 21140 13920 21146 13932
rect 21140 13892 21588 13920
rect 21140 13880 21146 13892
rect 19352 13824 20300 13852
rect 16868 13793 16896 13824
rect 20806 13812 20812 13864
rect 20864 13812 20870 13864
rect 21266 13812 21272 13864
rect 21324 13852 21330 13864
rect 21560 13852 21588 13892
rect 21726 13880 21732 13932
rect 21784 13920 21790 13932
rect 22020 13929 22048 13960
rect 21821 13923 21879 13929
rect 21821 13920 21833 13923
rect 21784 13892 21833 13920
rect 21784 13880 21790 13892
rect 21821 13889 21833 13892
rect 21867 13889 21879 13923
rect 21821 13883 21879 13889
rect 22005 13923 22063 13929
rect 22005 13889 22017 13923
rect 22051 13889 22063 13923
rect 22005 13883 22063 13889
rect 22097 13923 22155 13929
rect 22097 13889 22109 13923
rect 22143 13920 22155 13923
rect 23290 13920 23296 13932
rect 22143 13892 23296 13920
rect 22143 13889 22155 13892
rect 22097 13883 22155 13889
rect 23290 13880 23296 13892
rect 23348 13880 23354 13932
rect 24964 13929 24992 14028
rect 26418 14016 26424 14028
rect 26476 14016 26482 14068
rect 25041 13991 25099 13997
rect 25041 13957 25053 13991
rect 25087 13988 25099 13991
rect 27246 13988 27252 14000
rect 25087 13960 27252 13988
rect 25087 13957 25099 13960
rect 25041 13951 25099 13957
rect 27246 13948 27252 13960
rect 27304 13988 27310 14000
rect 27304 13960 27936 13988
rect 27304 13948 27310 13960
rect 24949 13923 25007 13929
rect 24949 13889 24961 13923
rect 24995 13889 25007 13923
rect 24949 13883 25007 13889
rect 25133 13923 25191 13929
rect 25133 13889 25145 13923
rect 25179 13889 25191 13923
rect 25133 13883 25191 13889
rect 25317 13923 25375 13929
rect 25317 13889 25329 13923
rect 25363 13920 25375 13923
rect 25774 13920 25780 13932
rect 25363 13892 25780 13920
rect 25363 13889 25375 13892
rect 25317 13883 25375 13889
rect 25148 13852 25176 13883
rect 25774 13880 25780 13892
rect 25832 13920 25838 13932
rect 25961 13923 26019 13929
rect 25961 13920 25973 13923
rect 25832 13892 25973 13920
rect 25832 13880 25838 13892
rect 25961 13889 25973 13892
rect 26007 13889 26019 13923
rect 25961 13883 26019 13889
rect 26326 13880 26332 13932
rect 26384 13880 26390 13932
rect 26694 13880 26700 13932
rect 26752 13880 26758 13932
rect 27908 13929 27936 13960
rect 27893 13923 27951 13929
rect 27893 13889 27905 13923
rect 27939 13889 27951 13923
rect 27893 13883 27951 13889
rect 28997 13923 29055 13929
rect 28997 13889 29009 13923
rect 29043 13920 29055 13923
rect 29457 13923 29515 13929
rect 29457 13920 29469 13923
rect 29043 13892 29469 13920
rect 29043 13889 29055 13892
rect 28997 13883 29055 13889
rect 29457 13889 29469 13892
rect 29503 13889 29515 13923
rect 29457 13883 29515 13889
rect 31202 13880 31208 13932
rect 31260 13880 31266 13932
rect 26712 13852 26740 13880
rect 21324 13824 21496 13852
rect 21560 13824 22094 13852
rect 21324 13812 21330 13824
rect 16853 13787 16911 13793
rect 16853 13784 16865 13787
rect 14976 13756 15608 13784
rect 15948 13756 16865 13784
rect 14976 13744 14982 13756
rect 15378 13676 15384 13728
rect 15436 13716 15442 13728
rect 15838 13716 15844 13728
rect 15436 13688 15844 13716
rect 15436 13676 15442 13688
rect 15838 13676 15844 13688
rect 15896 13716 15902 13728
rect 15948 13716 15976 13756
rect 16853 13753 16865 13756
rect 16899 13753 16911 13787
rect 16853 13747 16911 13753
rect 15896 13688 15976 13716
rect 15896 13676 15902 13688
rect 16022 13676 16028 13728
rect 16080 13716 16086 13728
rect 16117 13719 16175 13725
rect 16117 13716 16129 13719
rect 16080 13688 16129 13716
rect 16080 13676 16086 13688
rect 16117 13685 16129 13688
rect 16163 13685 16175 13719
rect 20824 13716 20852 13812
rect 21468 13793 21496 13824
rect 21453 13787 21511 13793
rect 21453 13753 21465 13787
rect 21499 13753 21511 13787
rect 22066 13784 22094 13824
rect 23400 13824 24808 13852
rect 25148 13824 26740 13852
rect 29089 13855 29147 13861
rect 22646 13784 22652 13796
rect 22066 13756 22652 13784
rect 21453 13747 21511 13753
rect 22646 13744 22652 13756
rect 22704 13744 22710 13796
rect 21726 13716 21732 13728
rect 20824 13688 21732 13716
rect 16117 13679 16175 13685
rect 21726 13676 21732 13688
rect 21784 13676 21790 13728
rect 22005 13719 22063 13725
rect 22005 13685 22017 13719
rect 22051 13716 22063 13719
rect 23400 13716 23428 13824
rect 24780 13793 24808 13824
rect 29089 13821 29101 13855
rect 29135 13821 29147 13855
rect 29089 13815 29147 13821
rect 29273 13855 29331 13861
rect 29273 13821 29285 13855
rect 29319 13852 29331 13855
rect 29638 13852 29644 13864
rect 29319 13824 29644 13852
rect 29319 13821 29331 13824
rect 29273 13815 29331 13821
rect 24765 13787 24823 13793
rect 24765 13753 24777 13787
rect 24811 13753 24823 13787
rect 29104 13784 29132 13815
rect 29638 13812 29644 13824
rect 29696 13812 29702 13864
rect 30098 13812 30104 13864
rect 30156 13812 30162 13864
rect 31478 13812 31484 13864
rect 31536 13812 31542 13864
rect 30006 13784 30012 13796
rect 24765 13747 24823 13753
rect 27448 13756 30012 13784
rect 27448 13728 27476 13756
rect 30006 13744 30012 13756
rect 30064 13744 30070 13796
rect 22051 13688 23428 13716
rect 22051 13685 22063 13688
rect 22005 13679 22063 13685
rect 25406 13676 25412 13728
rect 25464 13676 25470 13728
rect 26142 13676 26148 13728
rect 26200 13676 26206 13728
rect 27338 13676 27344 13728
rect 27396 13676 27402 13728
rect 27430 13676 27436 13728
rect 27488 13676 27494 13728
rect 27890 13676 27896 13728
rect 27948 13716 27954 13728
rect 28629 13719 28687 13725
rect 28629 13716 28641 13719
rect 27948 13688 28641 13716
rect 27948 13676 27954 13688
rect 28629 13685 28641 13688
rect 28675 13685 28687 13719
rect 28629 13679 28687 13685
rect 29362 13676 29368 13728
rect 29420 13716 29426 13728
rect 30116 13716 30144 13812
rect 29420 13688 30144 13716
rect 29420 13676 29426 13688
rect 1104 13626 31832 13648
rect 1104 13574 4182 13626
rect 4234 13574 4246 13626
rect 4298 13574 4310 13626
rect 4362 13574 4374 13626
rect 4426 13574 4438 13626
rect 4490 13574 4502 13626
rect 4554 13574 10182 13626
rect 10234 13574 10246 13626
rect 10298 13574 10310 13626
rect 10362 13574 10374 13626
rect 10426 13574 10438 13626
rect 10490 13574 10502 13626
rect 10554 13574 16182 13626
rect 16234 13574 16246 13626
rect 16298 13574 16310 13626
rect 16362 13574 16374 13626
rect 16426 13574 16438 13626
rect 16490 13574 16502 13626
rect 16554 13574 22182 13626
rect 22234 13574 22246 13626
rect 22298 13574 22310 13626
rect 22362 13574 22374 13626
rect 22426 13574 22438 13626
rect 22490 13574 22502 13626
rect 22554 13574 28182 13626
rect 28234 13574 28246 13626
rect 28298 13574 28310 13626
rect 28362 13574 28374 13626
rect 28426 13574 28438 13626
rect 28490 13574 28502 13626
rect 28554 13574 31832 13626
rect 1104 13552 31832 13574
rect 3234 13472 3240 13524
rect 3292 13512 3298 13524
rect 3789 13515 3847 13521
rect 3789 13512 3801 13515
rect 3292 13484 3801 13512
rect 3292 13472 3298 13484
rect 3789 13481 3801 13484
rect 3835 13481 3847 13515
rect 14093 13515 14151 13521
rect 14093 13512 14105 13515
rect 3789 13475 3847 13481
rect 12406 13484 14105 13512
rect 3786 13268 3792 13320
rect 3844 13308 3850 13320
rect 3973 13311 4031 13317
rect 3973 13308 3985 13311
rect 3844 13280 3985 13308
rect 3844 13268 3850 13280
rect 3973 13277 3985 13280
rect 4019 13277 4031 13311
rect 3973 13271 4031 13277
rect 12253 13311 12311 13317
rect 12253 13277 12265 13311
rect 12299 13308 12311 13311
rect 12406 13308 12434 13484
rect 14093 13481 14105 13484
rect 14139 13481 14151 13515
rect 14093 13475 14151 13481
rect 14826 13472 14832 13524
rect 14884 13512 14890 13524
rect 16206 13512 16212 13524
rect 14884 13484 16212 13512
rect 14884 13472 14890 13484
rect 16206 13472 16212 13484
rect 16264 13472 16270 13524
rect 18138 13472 18144 13524
rect 18196 13512 18202 13524
rect 19245 13515 19303 13521
rect 19245 13512 19257 13515
rect 18196 13484 19257 13512
rect 18196 13472 18202 13484
rect 19245 13481 19257 13484
rect 19291 13481 19303 13515
rect 19245 13475 19303 13481
rect 23290 13472 23296 13524
rect 23348 13512 23354 13524
rect 23348 13484 25728 13512
rect 23348 13472 23354 13484
rect 13909 13447 13967 13453
rect 13909 13413 13921 13447
rect 13955 13444 13967 13447
rect 13998 13444 14004 13456
rect 13955 13416 14004 13444
rect 13955 13413 13967 13416
rect 13909 13407 13967 13413
rect 13998 13404 14004 13416
rect 14056 13444 14062 13456
rect 22094 13444 22100 13456
rect 14056 13416 15516 13444
rect 14056 13404 14062 13416
rect 14090 13376 14096 13388
rect 13556 13348 14096 13376
rect 12299 13280 12434 13308
rect 12299 13277 12311 13280
rect 12253 13271 12311 13277
rect 12526 13268 12532 13320
rect 12584 13308 12590 13320
rect 13556 13308 13584 13348
rect 14090 13336 14096 13348
rect 14148 13336 14154 13388
rect 14550 13336 14556 13388
rect 14608 13336 14614 13388
rect 14642 13336 14648 13388
rect 14700 13336 14706 13388
rect 15488 13385 15516 13416
rect 19306 13416 22100 13444
rect 15473 13379 15531 13385
rect 15473 13345 15485 13379
rect 15519 13345 15531 13379
rect 19306 13376 19334 13416
rect 22094 13404 22100 13416
rect 22152 13404 22158 13456
rect 25700 13444 25728 13484
rect 25774 13472 25780 13524
rect 25832 13472 25838 13524
rect 25884 13484 26832 13512
rect 25884 13444 25912 13484
rect 25700 13416 25912 13444
rect 26804 13444 26832 13484
rect 27246 13472 27252 13524
rect 27304 13472 27310 13524
rect 27356 13484 29316 13512
rect 27356 13444 27384 13484
rect 26804 13416 27384 13444
rect 15473 13339 15531 13345
rect 15856 13348 19334 13376
rect 15856 13317 15884 13348
rect 19702 13336 19708 13388
rect 19760 13376 19766 13388
rect 19797 13379 19855 13385
rect 19797 13376 19809 13379
rect 19760 13348 19809 13376
rect 19760 13336 19766 13348
rect 19797 13345 19809 13348
rect 19843 13345 19855 13379
rect 19797 13339 19855 13345
rect 12584 13280 13584 13308
rect 15841 13311 15899 13317
rect 12584 13268 12590 13280
rect 15841 13277 15853 13311
rect 15887 13277 15899 13311
rect 15841 13271 15899 13277
rect 15933 13311 15991 13317
rect 15933 13277 15945 13311
rect 15979 13277 15991 13311
rect 15933 13271 15991 13277
rect 12774 13243 12832 13249
rect 12774 13240 12786 13243
rect 12452 13212 12786 13240
rect 12452 13181 12480 13212
rect 12774 13209 12786 13212
rect 12820 13209 12832 13243
rect 12774 13203 12832 13209
rect 14461 13243 14519 13249
rect 14461 13209 14473 13243
rect 14507 13240 14519 13243
rect 14921 13243 14979 13249
rect 14921 13240 14933 13243
rect 14507 13212 14933 13240
rect 14507 13209 14519 13212
rect 14461 13203 14519 13209
rect 14921 13209 14933 13212
rect 14967 13209 14979 13243
rect 15948 13240 15976 13271
rect 16022 13268 16028 13320
rect 16080 13268 16086 13320
rect 16114 13268 16120 13320
rect 16172 13268 16178 13320
rect 16206 13268 16212 13320
rect 16264 13308 16270 13320
rect 16301 13311 16359 13317
rect 16301 13308 16313 13311
rect 16264 13280 16313 13308
rect 16264 13268 16270 13280
rect 16301 13277 16313 13280
rect 16347 13277 16359 13311
rect 16301 13271 16359 13277
rect 16574 13268 16580 13320
rect 16632 13268 16638 13320
rect 24026 13268 24032 13320
rect 24084 13268 24090 13320
rect 24397 13311 24455 13317
rect 24397 13277 24409 13311
rect 24443 13308 24455 13311
rect 25869 13311 25927 13317
rect 25869 13308 25881 13311
rect 24443 13280 25881 13308
rect 24443 13277 24455 13280
rect 24397 13271 24455 13277
rect 25869 13277 25881 13280
rect 25915 13308 25927 13311
rect 26694 13308 26700 13320
rect 25915 13280 26700 13308
rect 25915 13277 25927 13280
rect 25869 13271 25927 13277
rect 26694 13268 26700 13280
rect 26752 13268 26758 13320
rect 27709 13311 27767 13317
rect 27709 13277 27721 13311
rect 27755 13308 27767 13311
rect 27890 13308 27896 13320
rect 27755 13280 27896 13308
rect 27755 13277 27767 13280
rect 27709 13271 27767 13277
rect 27890 13268 27896 13280
rect 27948 13268 27954 13320
rect 27985 13311 28043 13317
rect 27985 13277 27997 13311
rect 28031 13308 28043 13311
rect 28626 13308 28632 13320
rect 28031 13280 28632 13308
rect 28031 13277 28043 13280
rect 27985 13271 28043 13277
rect 28626 13268 28632 13280
rect 28684 13268 28690 13320
rect 26142 13249 26148 13252
rect 16761 13243 16819 13249
rect 16761 13240 16773 13243
rect 15948 13212 16773 13240
rect 14921 13203 14979 13209
rect 16761 13209 16773 13212
rect 16807 13209 16819 13243
rect 24642 13243 24700 13249
rect 24642 13240 24654 13243
rect 16761 13203 16819 13209
rect 24228 13212 24654 13240
rect 12437 13175 12495 13181
rect 12437 13141 12449 13175
rect 12483 13141 12495 13175
rect 12437 13135 12495 13141
rect 15654 13132 15660 13184
rect 15712 13132 15718 13184
rect 16022 13132 16028 13184
rect 16080 13172 16086 13184
rect 24228 13181 24256 13212
rect 24642 13209 24654 13212
rect 24688 13209 24700 13243
rect 26136 13240 26148 13249
rect 26103 13212 26148 13240
rect 24642 13203 24700 13209
rect 26136 13203 26148 13212
rect 26142 13200 26148 13203
rect 26200 13200 26206 13252
rect 28230 13243 28288 13249
rect 28230 13240 28242 13243
rect 27908 13212 28242 13240
rect 27908 13181 27936 13212
rect 28230 13209 28242 13212
rect 28276 13209 28288 13243
rect 28230 13203 28288 13209
rect 16393 13175 16451 13181
rect 16393 13172 16405 13175
rect 16080 13144 16405 13172
rect 16080 13132 16086 13144
rect 16393 13141 16405 13144
rect 16439 13141 16451 13175
rect 16393 13135 16451 13141
rect 24213 13175 24271 13181
rect 24213 13141 24225 13175
rect 24259 13141 24271 13175
rect 24213 13135 24271 13141
rect 27893 13175 27951 13181
rect 27893 13141 27905 13175
rect 27939 13141 27951 13175
rect 29288 13172 29316 13484
rect 29362 13472 29368 13524
rect 29420 13472 29426 13524
rect 29546 13472 29552 13524
rect 29604 13512 29610 13524
rect 29604 13484 30236 13512
rect 29604 13472 29610 13484
rect 29914 13404 29920 13456
rect 29972 13404 29978 13456
rect 29932 13376 29960 13404
rect 29702 13348 29960 13376
rect 29702 13317 29730 13348
rect 29687 13311 29745 13317
rect 29687 13277 29699 13311
rect 29733 13277 29745 13311
rect 30098 13308 30104 13320
rect 30059 13280 30104 13308
rect 29687 13271 29745 13277
rect 30098 13268 30104 13280
rect 30156 13268 30162 13320
rect 30208 13317 30236 13484
rect 30193 13311 30251 13317
rect 30193 13277 30205 13311
rect 30239 13277 30251 13311
rect 30193 13271 30251 13277
rect 29822 13200 29828 13252
rect 29880 13200 29886 13252
rect 29917 13243 29975 13249
rect 29917 13209 29929 13243
rect 29963 13240 29975 13243
rect 30650 13240 30656 13252
rect 29963 13212 30656 13240
rect 29963 13209 29975 13212
rect 29917 13203 29975 13209
rect 30650 13200 30656 13212
rect 30708 13200 30714 13252
rect 29549 13175 29607 13181
rect 29549 13172 29561 13175
rect 29288 13144 29561 13172
rect 27893 13135 27951 13141
rect 29549 13141 29561 13144
rect 29595 13141 29607 13175
rect 29549 13135 29607 13141
rect 29730 13132 29736 13184
rect 29788 13172 29794 13184
rect 30190 13172 30196 13184
rect 29788 13144 30196 13172
rect 29788 13132 29794 13144
rect 30190 13132 30196 13144
rect 30248 13132 30254 13184
rect 1104 13082 31832 13104
rect 1104 13030 4922 13082
rect 4974 13030 4986 13082
rect 5038 13030 5050 13082
rect 5102 13030 5114 13082
rect 5166 13030 5178 13082
rect 5230 13030 5242 13082
rect 5294 13030 10922 13082
rect 10974 13030 10986 13082
rect 11038 13030 11050 13082
rect 11102 13030 11114 13082
rect 11166 13030 11178 13082
rect 11230 13030 11242 13082
rect 11294 13030 16922 13082
rect 16974 13030 16986 13082
rect 17038 13030 17050 13082
rect 17102 13030 17114 13082
rect 17166 13030 17178 13082
rect 17230 13030 17242 13082
rect 17294 13030 22922 13082
rect 22974 13030 22986 13082
rect 23038 13030 23050 13082
rect 23102 13030 23114 13082
rect 23166 13030 23178 13082
rect 23230 13030 23242 13082
rect 23294 13030 28922 13082
rect 28974 13030 28986 13082
rect 29038 13030 29050 13082
rect 29102 13030 29114 13082
rect 29166 13030 29178 13082
rect 29230 13030 29242 13082
rect 29294 13030 31832 13082
rect 1104 13008 31832 13030
rect 9766 12968 9772 12980
rect 2746 12940 9772 12968
rect 1765 12903 1823 12909
rect 1765 12869 1777 12903
rect 1811 12900 1823 12903
rect 2746 12900 2774 12940
rect 9766 12928 9772 12940
rect 9824 12968 9830 12980
rect 10413 12971 10471 12977
rect 10413 12968 10425 12971
rect 9824 12940 10425 12968
rect 9824 12928 9830 12940
rect 10413 12937 10425 12940
rect 10459 12937 10471 12971
rect 10413 12931 10471 12937
rect 13998 12928 14004 12980
rect 14056 12928 14062 12980
rect 14277 12971 14335 12977
rect 14277 12937 14289 12971
rect 14323 12968 14335 12971
rect 15930 12968 15936 12980
rect 14323 12940 15936 12968
rect 14323 12937 14335 12940
rect 14277 12931 14335 12937
rect 15930 12928 15936 12940
rect 15988 12928 15994 12980
rect 22646 12928 22652 12980
rect 22704 12928 22710 12980
rect 24026 12928 24032 12980
rect 24084 12968 24090 12980
rect 24489 12971 24547 12977
rect 24489 12968 24501 12971
rect 24084 12940 24501 12968
rect 24084 12928 24090 12940
rect 24489 12937 24501 12940
rect 24535 12937 24547 12971
rect 24489 12931 24547 12937
rect 24857 12971 24915 12977
rect 24857 12937 24869 12971
rect 24903 12968 24915 12971
rect 25406 12968 25412 12980
rect 24903 12940 25412 12968
rect 24903 12937 24915 12940
rect 24857 12931 24915 12937
rect 25406 12928 25412 12940
rect 25464 12928 25470 12980
rect 26326 12928 26332 12980
rect 26384 12968 26390 12980
rect 26973 12971 27031 12977
rect 26973 12968 26985 12971
rect 26384 12940 26985 12968
rect 26384 12928 26390 12940
rect 26973 12937 26985 12940
rect 27019 12937 27031 12971
rect 26973 12931 27031 12937
rect 27338 12928 27344 12980
rect 27396 12928 27402 12980
rect 28537 12971 28595 12977
rect 28537 12937 28549 12971
rect 28583 12968 28595 12971
rect 28583 12940 28764 12968
rect 28583 12937 28595 12940
rect 28537 12931 28595 12937
rect 9030 12900 9036 12912
rect 1811 12872 2774 12900
rect 8680 12872 9036 12900
rect 1811 12869 1823 12872
rect 1765 12863 1823 12869
rect 8294 12792 8300 12844
rect 8352 12832 8358 12844
rect 8680 12841 8708 12872
rect 9030 12860 9036 12872
rect 9088 12860 9094 12912
rect 10597 12903 10655 12909
rect 10597 12900 10609 12903
rect 10166 12872 10609 12900
rect 10597 12869 10609 12872
rect 10643 12869 10655 12903
rect 10597 12863 10655 12869
rect 12894 12860 12900 12912
rect 12952 12900 12958 12912
rect 12989 12903 13047 12909
rect 12989 12900 13001 12903
rect 12952 12872 13001 12900
rect 12952 12860 12958 12872
rect 12989 12869 13001 12872
rect 13035 12900 13047 12903
rect 13262 12900 13268 12912
rect 13035 12872 13268 12900
rect 13035 12869 13047 12872
rect 12989 12863 13047 12869
rect 13262 12860 13268 12872
rect 13320 12860 13326 12912
rect 13446 12860 13452 12912
rect 13504 12900 13510 12912
rect 13504 12872 13768 12900
rect 13504 12860 13510 12872
rect 8665 12835 8723 12841
rect 8665 12832 8677 12835
rect 8352 12804 8677 12832
rect 8352 12792 8358 12804
rect 8665 12801 8677 12804
rect 8711 12801 8723 12835
rect 8665 12795 8723 12801
rect 10689 12835 10747 12841
rect 10689 12801 10701 12835
rect 10735 12801 10747 12835
rect 10689 12795 10747 12801
rect 8938 12724 8944 12776
rect 8996 12724 9002 12776
rect 9674 12724 9680 12776
rect 9732 12764 9738 12776
rect 10704 12764 10732 12795
rect 12618 12792 12624 12844
rect 12676 12792 12682 12844
rect 12802 12792 12808 12844
rect 12860 12792 12866 12844
rect 13078 12792 13084 12844
rect 13136 12792 13142 12844
rect 13740 12841 13768 12872
rect 13814 12860 13820 12912
rect 13872 12900 13878 12912
rect 13909 12903 13967 12909
rect 13909 12900 13921 12903
rect 13872 12872 13921 12900
rect 13872 12860 13878 12872
rect 13909 12869 13921 12872
rect 13955 12869 13967 12903
rect 13909 12863 13967 12869
rect 14016 12841 14044 12928
rect 22664 12900 22692 12928
rect 24949 12903 25007 12909
rect 24949 12900 24961 12903
rect 22664 12872 24961 12900
rect 24949 12869 24961 12872
rect 24995 12900 25007 12903
rect 24995 12872 26648 12900
rect 24995 12869 25007 12872
rect 24949 12863 25007 12869
rect 14182 12841 14188 12844
rect 13173 12835 13231 12841
rect 13173 12801 13185 12835
rect 13219 12801 13231 12835
rect 13633 12835 13691 12841
rect 13633 12832 13645 12835
rect 13173 12795 13231 12801
rect 13372 12804 13645 12832
rect 9732 12736 10732 12764
rect 12636 12764 12664 12792
rect 13188 12764 13216 12795
rect 12636 12736 13216 12764
rect 9732 12724 9738 12736
rect 10060 12708 10088 12736
rect 10042 12656 10048 12708
rect 10100 12656 10106 12708
rect 1486 12588 1492 12640
rect 1544 12588 1550 12640
rect 13188 12628 13216 12736
rect 13372 12705 13400 12804
rect 13633 12801 13645 12804
rect 13679 12801 13691 12835
rect 13633 12795 13691 12801
rect 13726 12835 13784 12841
rect 13726 12801 13738 12835
rect 13772 12801 13784 12835
rect 13726 12795 13784 12801
rect 14001 12835 14059 12841
rect 14001 12801 14013 12835
rect 14047 12801 14059 12835
rect 14001 12795 14059 12801
rect 14139 12835 14188 12841
rect 14139 12801 14151 12835
rect 14185 12801 14188 12835
rect 14139 12795 14188 12801
rect 14182 12792 14188 12795
rect 14240 12832 14246 12844
rect 14366 12832 14372 12844
rect 14240 12804 14372 12832
rect 14240 12792 14246 12804
rect 14366 12792 14372 12804
rect 14424 12792 14430 12844
rect 20530 12792 20536 12844
rect 20588 12792 20594 12844
rect 22189 12835 22247 12841
rect 22189 12801 22201 12835
rect 22235 12832 22247 12835
rect 22922 12832 22928 12844
rect 22235 12804 22928 12832
rect 22235 12801 22247 12804
rect 22189 12795 22247 12801
rect 22922 12792 22928 12804
rect 22980 12792 22986 12844
rect 25406 12792 25412 12844
rect 25464 12832 25470 12844
rect 25869 12835 25927 12841
rect 25869 12832 25881 12835
rect 25464 12804 25881 12832
rect 25464 12792 25470 12804
rect 25869 12801 25881 12804
rect 25915 12801 25927 12835
rect 26620 12832 26648 12872
rect 26694 12860 26700 12912
rect 26752 12900 26758 12912
rect 28736 12900 28764 12940
rect 29362 12928 29368 12980
rect 29420 12968 29426 12980
rect 29546 12968 29552 12980
rect 29420 12940 29552 12968
rect 29420 12928 29426 12940
rect 29546 12928 29552 12940
rect 29604 12928 29610 12980
rect 29822 12928 29828 12980
rect 29880 12968 29886 12980
rect 30009 12971 30067 12977
rect 30009 12968 30021 12971
rect 29880 12940 30021 12968
rect 29880 12928 29886 12940
rect 30009 12937 30021 12940
rect 30055 12937 30067 12971
rect 30009 12931 30067 12937
rect 28874 12903 28932 12909
rect 28874 12900 28886 12903
rect 26752 12872 28672 12900
rect 28736 12872 28886 12900
rect 26752 12860 26758 12872
rect 28644 12844 28672 12872
rect 28874 12869 28886 12872
rect 28920 12869 28932 12903
rect 28874 12863 28932 12869
rect 27430 12832 27436 12844
rect 26620 12804 27436 12832
rect 25869 12795 25927 12801
rect 27430 12792 27436 12804
rect 27488 12792 27494 12844
rect 28353 12835 28411 12841
rect 28353 12801 28365 12835
rect 28399 12832 28411 12835
rect 28399 12804 28488 12832
rect 28399 12801 28411 12804
rect 28353 12795 28411 12801
rect 21361 12767 21419 12773
rect 21361 12733 21373 12767
rect 21407 12764 21419 12767
rect 21450 12764 21456 12776
rect 21407 12736 21456 12764
rect 21407 12733 21419 12736
rect 21361 12727 21419 12733
rect 21450 12724 21456 12736
rect 21508 12724 21514 12776
rect 23842 12724 23848 12776
rect 23900 12724 23906 12776
rect 25133 12767 25191 12773
rect 25133 12733 25145 12767
rect 25179 12764 25191 12767
rect 25222 12764 25228 12776
rect 25179 12736 25228 12764
rect 25179 12733 25191 12736
rect 25133 12727 25191 12733
rect 25222 12724 25228 12736
rect 25280 12724 25286 12776
rect 27062 12724 27068 12776
rect 27120 12764 27126 12776
rect 27522 12764 27528 12776
rect 27120 12736 27528 12764
rect 27120 12724 27126 12736
rect 27522 12724 27528 12736
rect 27580 12724 27586 12776
rect 13357 12699 13415 12705
rect 13357 12665 13369 12699
rect 13403 12665 13415 12699
rect 13357 12659 13415 12665
rect 13538 12628 13544 12640
rect 13188 12600 13544 12628
rect 13538 12588 13544 12600
rect 13596 12588 13602 12640
rect 22005 12631 22063 12637
rect 22005 12597 22017 12631
rect 22051 12628 22063 12631
rect 22094 12628 22100 12640
rect 22051 12600 22100 12628
rect 22051 12597 22063 12600
rect 22005 12591 22063 12597
rect 22094 12588 22100 12600
rect 22152 12588 22158 12640
rect 23290 12588 23296 12640
rect 23348 12588 23354 12640
rect 28460 12628 28488 12804
rect 28626 12792 28632 12844
rect 28684 12792 28690 12844
rect 30024 12832 30052 12931
rect 30653 12835 30711 12841
rect 30653 12832 30665 12835
rect 30024 12804 30665 12832
rect 30653 12801 30665 12804
rect 30699 12801 30711 12835
rect 30653 12795 30711 12801
rect 29546 12628 29552 12640
rect 28460 12600 29552 12628
rect 29546 12588 29552 12600
rect 29604 12588 29610 12640
rect 30098 12588 30104 12640
rect 30156 12588 30162 12640
rect 1104 12538 31832 12560
rect 1104 12486 4182 12538
rect 4234 12486 4246 12538
rect 4298 12486 4310 12538
rect 4362 12486 4374 12538
rect 4426 12486 4438 12538
rect 4490 12486 4502 12538
rect 4554 12486 10182 12538
rect 10234 12486 10246 12538
rect 10298 12486 10310 12538
rect 10362 12486 10374 12538
rect 10426 12486 10438 12538
rect 10490 12486 10502 12538
rect 10554 12486 16182 12538
rect 16234 12486 16246 12538
rect 16298 12486 16310 12538
rect 16362 12486 16374 12538
rect 16426 12486 16438 12538
rect 16490 12486 16502 12538
rect 16554 12486 22182 12538
rect 22234 12486 22246 12538
rect 22298 12486 22310 12538
rect 22362 12486 22374 12538
rect 22426 12486 22438 12538
rect 22490 12486 22502 12538
rect 22554 12486 28182 12538
rect 28234 12486 28246 12538
rect 28298 12486 28310 12538
rect 28362 12486 28374 12538
rect 28426 12486 28438 12538
rect 28490 12486 28502 12538
rect 28554 12486 31832 12538
rect 1104 12464 31832 12486
rect 8938 12384 8944 12436
rect 8996 12424 9002 12436
rect 9125 12427 9183 12433
rect 9125 12424 9137 12427
rect 8996 12396 9137 12424
rect 8996 12384 9002 12396
rect 9125 12393 9137 12396
rect 9171 12393 9183 12427
rect 9125 12387 9183 12393
rect 22922 12384 22928 12436
rect 22980 12384 22986 12436
rect 29546 12384 29552 12436
rect 29604 12384 29610 12436
rect 5442 12316 5448 12368
rect 5500 12356 5506 12368
rect 5500 12328 7972 12356
rect 5500 12316 5506 12328
rect 4154 12248 4160 12300
rect 4212 12288 4218 12300
rect 4706 12288 4712 12300
rect 4212 12260 4712 12288
rect 4212 12248 4218 12260
rect 4706 12248 4712 12260
rect 4764 12288 4770 12300
rect 6089 12291 6147 12297
rect 6089 12288 6101 12291
rect 4764 12260 6101 12288
rect 4764 12248 4770 12260
rect 6089 12257 6101 12260
rect 6135 12257 6147 12291
rect 6089 12251 6147 12257
rect 6273 12291 6331 12297
rect 6273 12257 6285 12291
rect 6319 12288 6331 12291
rect 7190 12288 7196 12300
rect 6319 12260 7196 12288
rect 6319 12257 6331 12260
rect 6273 12251 6331 12257
rect 7190 12248 7196 12260
rect 7248 12248 7254 12300
rect 4798 12220 4804 12232
rect 3988 12192 4804 12220
rect 3988 12096 4016 12192
rect 4798 12180 4804 12192
rect 4856 12220 4862 12232
rect 4893 12223 4951 12229
rect 4893 12220 4905 12223
rect 4856 12192 4905 12220
rect 4856 12180 4862 12192
rect 4893 12189 4905 12192
rect 4939 12189 4951 12223
rect 4893 12183 4951 12189
rect 5169 12223 5227 12229
rect 5169 12189 5181 12223
rect 5215 12189 5227 12223
rect 5169 12183 5227 12189
rect 4706 12112 4712 12164
rect 4764 12152 4770 12164
rect 5184 12152 5212 12183
rect 7006 12180 7012 12232
rect 7064 12180 7070 12232
rect 7098 12152 7104 12164
rect 4764 12124 5212 12152
rect 6748 12124 7104 12152
rect 4764 12112 4770 12124
rect 3970 12044 3976 12096
rect 4028 12044 4034 12096
rect 4246 12044 4252 12096
rect 4304 12044 4310 12096
rect 4430 12044 4436 12096
rect 4488 12084 4494 12096
rect 4985 12087 5043 12093
rect 4985 12084 4997 12087
rect 4488 12056 4997 12084
rect 4488 12044 4494 12056
rect 4985 12053 4997 12056
rect 5031 12053 5043 12087
rect 4985 12047 5043 12053
rect 6362 12044 6368 12096
rect 6420 12044 6426 12096
rect 6748 12093 6776 12124
rect 7098 12112 7104 12124
rect 7156 12112 7162 12164
rect 7944 12096 7972 12328
rect 9674 12316 9680 12368
rect 9732 12356 9738 12368
rect 10042 12356 10048 12368
rect 9732 12328 10048 12356
rect 9732 12316 9738 12328
rect 10042 12316 10048 12328
rect 10100 12316 10106 12368
rect 9950 12248 9956 12300
rect 10008 12248 10014 12300
rect 15286 12248 15292 12300
rect 15344 12288 15350 12300
rect 15562 12288 15568 12300
rect 15344 12260 15568 12288
rect 15344 12248 15350 12260
rect 15562 12248 15568 12260
rect 15620 12288 15626 12300
rect 15657 12291 15715 12297
rect 15657 12288 15669 12291
rect 15620 12260 15669 12288
rect 15620 12248 15626 12260
rect 15657 12257 15669 12260
rect 15703 12257 15715 12291
rect 15657 12251 15715 12257
rect 15838 12248 15844 12300
rect 15896 12248 15902 12300
rect 19889 12291 19947 12297
rect 19889 12257 19901 12291
rect 19935 12288 19947 12291
rect 19935 12260 21312 12288
rect 19935 12257 19947 12260
rect 19889 12251 19947 12257
rect 8018 12180 8024 12232
rect 8076 12180 8082 12232
rect 8662 12180 8668 12232
rect 8720 12180 8726 12232
rect 9309 12223 9367 12229
rect 9309 12189 9321 12223
rect 9355 12220 9367 12223
rect 9355 12192 9444 12220
rect 9355 12189 9367 12192
rect 9309 12183 9367 12189
rect 6733 12087 6791 12093
rect 6733 12053 6745 12087
rect 6779 12053 6791 12087
rect 6733 12047 6791 12053
rect 6822 12044 6828 12096
rect 6880 12044 6886 12096
rect 6914 12044 6920 12096
rect 6972 12084 6978 12096
rect 7377 12087 7435 12093
rect 7377 12084 7389 12087
rect 6972 12056 7389 12084
rect 6972 12044 6978 12056
rect 7377 12053 7389 12056
rect 7423 12053 7435 12087
rect 7377 12047 7435 12053
rect 7926 12044 7932 12096
rect 7984 12044 7990 12096
rect 8478 12044 8484 12096
rect 8536 12044 8542 12096
rect 9416 12093 9444 12192
rect 9766 12180 9772 12232
rect 9824 12180 9830 12232
rect 16114 12180 16120 12232
rect 16172 12220 16178 12232
rect 16945 12223 17003 12229
rect 16945 12220 16957 12223
rect 16172 12192 16957 12220
rect 16172 12180 16178 12192
rect 16945 12189 16957 12192
rect 16991 12189 17003 12223
rect 16945 12183 17003 12189
rect 20809 12223 20867 12229
rect 20809 12189 20821 12223
rect 20855 12220 20867 12223
rect 21177 12223 21235 12229
rect 20855 12192 21128 12220
rect 20855 12189 20867 12192
rect 20809 12183 20867 12189
rect 15933 12155 15991 12161
rect 15933 12121 15945 12155
rect 15979 12152 15991 12155
rect 16393 12155 16451 12161
rect 16393 12152 16405 12155
rect 15979 12124 16405 12152
rect 15979 12121 15991 12124
rect 15933 12115 15991 12121
rect 16393 12121 16405 12124
rect 16439 12121 16451 12155
rect 16393 12115 16451 12121
rect 19613 12155 19671 12161
rect 19613 12121 19625 12155
rect 19659 12152 19671 12155
rect 20165 12155 20223 12161
rect 20165 12152 20177 12155
rect 19659 12124 20177 12152
rect 19659 12121 19671 12124
rect 19613 12115 19671 12121
rect 20165 12121 20177 12124
rect 20211 12121 20223 12155
rect 20165 12115 20223 12121
rect 21100 12096 21128 12192
rect 21177 12189 21189 12223
rect 21223 12189 21235 12223
rect 21284 12220 21312 12260
rect 21450 12248 21456 12300
rect 21508 12248 21514 12300
rect 23569 12291 23627 12297
rect 23569 12288 23581 12291
rect 23216 12260 23581 12288
rect 23216 12220 23244 12260
rect 23569 12257 23581 12260
rect 23615 12288 23627 12291
rect 27522 12288 27528 12300
rect 23615 12260 27528 12288
rect 23615 12257 23627 12260
rect 23569 12251 23627 12257
rect 27522 12248 27528 12260
rect 27580 12248 27586 12300
rect 30006 12248 30012 12300
rect 30064 12248 30070 12300
rect 30190 12248 30196 12300
rect 30248 12248 30254 12300
rect 21284 12192 23244 12220
rect 21177 12183 21235 12189
rect 21192 12152 21220 12183
rect 23290 12180 23296 12232
rect 23348 12180 23354 12232
rect 21266 12152 21272 12164
rect 21192 12124 21272 12152
rect 21266 12112 21272 12124
rect 21324 12112 21330 12164
rect 21698 12155 21756 12161
rect 21698 12152 21710 12155
rect 21376 12124 21710 12152
rect 9401 12087 9459 12093
rect 9401 12053 9413 12087
rect 9447 12053 9459 12087
rect 9401 12047 9459 12053
rect 9861 12087 9919 12093
rect 9861 12053 9873 12087
rect 9907 12084 9919 12087
rect 10042 12084 10048 12096
rect 9907 12056 10048 12084
rect 9907 12053 9919 12056
rect 9861 12047 9919 12053
rect 10042 12044 10048 12056
rect 10100 12044 10106 12096
rect 16022 12044 16028 12096
rect 16080 12084 16086 12096
rect 16301 12087 16359 12093
rect 16301 12084 16313 12087
rect 16080 12056 16313 12084
rect 16080 12044 16086 12056
rect 16301 12053 16313 12056
rect 16347 12053 16359 12087
rect 16301 12047 16359 12053
rect 19242 12044 19248 12096
rect 19300 12044 19306 12096
rect 19702 12044 19708 12096
rect 19760 12044 19766 12096
rect 21082 12044 21088 12096
rect 21140 12044 21146 12096
rect 21376 12093 21404 12124
rect 21698 12121 21710 12124
rect 21744 12121 21756 12155
rect 21698 12115 21756 12121
rect 25406 12112 25412 12164
rect 25464 12112 25470 12164
rect 26050 12112 26056 12164
rect 26108 12152 26114 12164
rect 26145 12155 26203 12161
rect 26145 12152 26157 12155
rect 26108 12124 26157 12152
rect 26108 12112 26114 12124
rect 26145 12121 26157 12124
rect 26191 12121 26203 12155
rect 26145 12115 26203 12121
rect 29917 12155 29975 12161
rect 29917 12121 29929 12155
rect 29963 12152 29975 12155
rect 30098 12152 30104 12164
rect 29963 12124 30104 12152
rect 29963 12121 29975 12124
rect 29917 12115 29975 12121
rect 30098 12112 30104 12124
rect 30156 12112 30162 12164
rect 21361 12087 21419 12093
rect 21361 12053 21373 12087
rect 21407 12053 21419 12087
rect 21361 12047 21419 12053
rect 22830 12044 22836 12096
rect 22888 12044 22894 12096
rect 23385 12087 23443 12093
rect 23385 12053 23397 12087
rect 23431 12084 23443 12087
rect 24670 12084 24676 12096
rect 23431 12056 24676 12084
rect 23431 12053 23443 12056
rect 23385 12047 23443 12053
rect 24670 12044 24676 12056
rect 24728 12044 24734 12096
rect 1104 11994 31832 12016
rect 1104 11942 4922 11994
rect 4974 11942 4986 11994
rect 5038 11942 5050 11994
rect 5102 11942 5114 11994
rect 5166 11942 5178 11994
rect 5230 11942 5242 11994
rect 5294 11942 10922 11994
rect 10974 11942 10986 11994
rect 11038 11942 11050 11994
rect 11102 11942 11114 11994
rect 11166 11942 11178 11994
rect 11230 11942 11242 11994
rect 11294 11942 16922 11994
rect 16974 11942 16986 11994
rect 17038 11942 17050 11994
rect 17102 11942 17114 11994
rect 17166 11942 17178 11994
rect 17230 11942 17242 11994
rect 17294 11942 22922 11994
rect 22974 11942 22986 11994
rect 23038 11942 23050 11994
rect 23102 11942 23114 11994
rect 23166 11942 23178 11994
rect 23230 11942 23242 11994
rect 23294 11942 28922 11994
rect 28974 11942 28986 11994
rect 29038 11942 29050 11994
rect 29102 11942 29114 11994
rect 29166 11942 29178 11994
rect 29230 11942 29242 11994
rect 29294 11942 31832 11994
rect 1104 11920 31832 11942
rect 3970 11840 3976 11892
rect 4028 11840 4034 11892
rect 4246 11840 4252 11892
rect 4304 11880 4310 11892
rect 4433 11883 4491 11889
rect 4433 11880 4445 11883
rect 4304 11852 4445 11880
rect 4304 11840 4310 11852
rect 4433 11849 4445 11852
rect 4479 11849 4491 11883
rect 4433 11843 4491 11849
rect 4706 11840 4712 11892
rect 4764 11880 4770 11892
rect 4801 11883 4859 11889
rect 4801 11880 4813 11883
rect 4764 11852 4813 11880
rect 4764 11840 4770 11852
rect 4801 11849 4813 11852
rect 4847 11849 4859 11883
rect 4801 11843 4859 11849
rect 5074 11840 5080 11892
rect 5132 11880 5138 11892
rect 5442 11880 5448 11892
rect 5132 11852 5448 11880
rect 5132 11840 5138 11852
rect 5442 11840 5448 11852
rect 5500 11840 5506 11892
rect 6181 11883 6239 11889
rect 6181 11849 6193 11883
rect 6227 11880 6239 11883
rect 6362 11880 6368 11892
rect 6227 11852 6368 11880
rect 6227 11849 6239 11852
rect 6181 11843 6239 11849
rect 6362 11840 6368 11852
rect 6420 11840 6426 11892
rect 6822 11840 6828 11892
rect 6880 11840 6886 11892
rect 7745 11883 7803 11889
rect 7745 11849 7757 11883
rect 7791 11880 7803 11883
rect 8018 11880 8024 11892
rect 7791 11852 8024 11880
rect 7791 11849 7803 11852
rect 7745 11843 7803 11849
rect 8018 11840 8024 11852
rect 8076 11880 8082 11892
rect 8076 11852 8156 11880
rect 8076 11840 8082 11852
rect 6632 11815 6690 11821
rect 2608 11784 6408 11812
rect 2608 11756 2636 11784
rect 6380 11756 6408 11784
rect 6632 11781 6644 11815
rect 6678 11812 6690 11815
rect 6840 11812 6868 11840
rect 8128 11821 8156 11852
rect 16114 11840 16120 11892
rect 16172 11880 16178 11892
rect 16485 11883 16543 11889
rect 16485 11880 16497 11883
rect 16172 11852 16497 11880
rect 16172 11840 16178 11852
rect 16485 11849 16497 11852
rect 16531 11849 16543 11883
rect 16485 11843 16543 11849
rect 23201 11883 23259 11889
rect 23201 11849 23213 11883
rect 23247 11880 23259 11883
rect 23842 11880 23848 11892
rect 23247 11852 23848 11880
rect 23247 11849 23259 11852
rect 23201 11843 23259 11849
rect 23842 11840 23848 11852
rect 23900 11840 23906 11892
rect 6678 11784 6868 11812
rect 8113 11815 8171 11821
rect 6678 11781 6690 11784
rect 6632 11775 6690 11781
rect 8113 11781 8125 11815
rect 8159 11781 8171 11815
rect 8113 11775 8171 11781
rect 19168 11784 19840 11812
rect 2590 11704 2596 11756
rect 2648 11704 2654 11756
rect 2860 11747 2918 11753
rect 2860 11713 2872 11747
rect 2906 11744 2918 11747
rect 4430 11744 4436 11756
rect 2906 11716 4436 11744
rect 2906 11713 2918 11716
rect 2860 11707 2918 11713
rect 4430 11704 4436 11716
rect 4488 11704 4494 11756
rect 4798 11704 4804 11756
rect 4856 11744 4862 11756
rect 4893 11747 4951 11753
rect 4893 11744 4905 11747
rect 4856 11716 4905 11744
rect 4856 11704 4862 11716
rect 4893 11713 4905 11716
rect 4939 11713 4951 11747
rect 4893 11707 4951 11713
rect 5074 11704 5080 11756
rect 5132 11704 5138 11756
rect 5166 11704 5172 11756
rect 5224 11704 5230 11756
rect 5261 11747 5319 11753
rect 5261 11713 5273 11747
rect 5307 11744 5319 11747
rect 5350 11744 5356 11756
rect 5307 11716 5356 11744
rect 5307 11713 5319 11716
rect 5261 11707 5319 11713
rect 5350 11704 5356 11716
rect 5408 11744 5414 11756
rect 6178 11744 6184 11756
rect 5408 11716 6184 11744
rect 5408 11704 5414 11716
rect 6178 11704 6184 11716
rect 6236 11704 6242 11756
rect 6362 11704 6368 11756
rect 6420 11704 6426 11756
rect 7837 11747 7895 11753
rect 7837 11744 7849 11747
rect 6472 11716 7849 11744
rect 3694 11636 3700 11688
rect 3752 11636 3758 11688
rect 4154 11636 4160 11688
rect 4212 11636 4218 11688
rect 4341 11679 4399 11685
rect 4341 11645 4353 11679
rect 4387 11645 4399 11679
rect 4341 11639 4399 11645
rect 3712 11608 3740 11636
rect 4356 11608 4384 11639
rect 5626 11636 5632 11688
rect 5684 11676 5690 11688
rect 6472 11676 6500 11716
rect 7837 11713 7849 11716
rect 7883 11713 7895 11747
rect 7837 11707 7895 11713
rect 7926 11704 7932 11756
rect 7984 11744 7990 11756
rect 8021 11747 8079 11753
rect 8021 11744 8033 11747
rect 7984 11716 8033 11744
rect 7984 11704 7990 11716
rect 8021 11713 8033 11716
rect 8067 11713 8079 11747
rect 8021 11707 8079 11713
rect 8205 11747 8263 11753
rect 8205 11713 8217 11747
rect 8251 11713 8263 11747
rect 8205 11707 8263 11713
rect 9401 11747 9459 11753
rect 9401 11713 9413 11747
rect 9447 11744 9459 11747
rect 9858 11744 9864 11756
rect 9447 11716 9864 11744
rect 9447 11713 9459 11716
rect 9401 11707 9459 11713
rect 5684 11648 6500 11676
rect 5684 11636 5690 11648
rect 7374 11636 7380 11688
rect 7432 11676 7438 11688
rect 8220 11676 8248 11707
rect 9858 11704 9864 11716
rect 9916 11704 9922 11756
rect 13725 11747 13783 11753
rect 13725 11713 13737 11747
rect 13771 11744 13783 11747
rect 14182 11744 14188 11756
rect 13771 11716 14188 11744
rect 13771 11713 13783 11716
rect 13725 11707 13783 11713
rect 14182 11704 14188 11716
rect 14240 11704 14246 11756
rect 15372 11747 15430 11753
rect 15372 11713 15384 11747
rect 15418 11744 15430 11747
rect 15930 11744 15936 11756
rect 15418 11716 15936 11744
rect 15418 11713 15430 11716
rect 15372 11707 15430 11713
rect 15930 11704 15936 11716
rect 15988 11704 15994 11756
rect 17954 11753 17960 11756
rect 17948 11707 17960 11753
rect 17954 11704 17960 11707
rect 18012 11704 18018 11756
rect 7432 11648 8248 11676
rect 8665 11679 8723 11685
rect 7432 11636 7438 11648
rect 8665 11645 8677 11679
rect 8711 11676 8723 11679
rect 8938 11676 8944 11688
rect 8711 11648 8944 11676
rect 8711 11645 8723 11648
rect 8665 11639 8723 11645
rect 8938 11636 8944 11648
rect 8996 11636 9002 11688
rect 13998 11636 14004 11688
rect 14056 11676 14062 11688
rect 19168 11685 19196 11784
rect 19426 11753 19432 11756
rect 19420 11707 19432 11753
rect 19426 11704 19432 11707
rect 19484 11704 19490 11756
rect 19812 11744 19840 11784
rect 20714 11772 20720 11824
rect 20772 11812 20778 11824
rect 21545 11815 21603 11821
rect 21545 11812 21557 11815
rect 20772 11784 21557 11812
rect 20772 11772 20778 11784
rect 21545 11781 21557 11784
rect 21591 11812 21603 11815
rect 21634 11812 21640 11824
rect 21591 11784 21640 11812
rect 21591 11781 21603 11784
rect 21545 11775 21603 11781
rect 21634 11772 21640 11784
rect 21692 11772 21698 11824
rect 22094 11821 22100 11824
rect 22088 11775 22100 11821
rect 22152 11812 22158 11824
rect 22152 11784 22188 11812
rect 22094 11772 22100 11775
rect 22152 11772 22158 11784
rect 22278 11772 22284 11824
rect 22336 11812 22342 11824
rect 23293 11815 23351 11821
rect 23293 11812 23305 11815
rect 22336 11784 23305 11812
rect 22336 11772 22342 11784
rect 23293 11781 23305 11784
rect 23339 11781 23351 11815
rect 23293 11775 23351 11781
rect 26510 11772 26516 11824
rect 26568 11772 26574 11824
rect 20809 11747 20867 11753
rect 20809 11744 20821 11747
rect 19812 11716 20821 11744
rect 20809 11713 20821 11716
rect 20855 11744 20867 11747
rect 21821 11747 21879 11753
rect 21821 11744 21833 11747
rect 20855 11716 21833 11744
rect 20855 11713 20867 11716
rect 20809 11707 20867 11713
rect 21821 11713 21833 11716
rect 21867 11713 21879 11747
rect 21821 11707 21879 11713
rect 22830 11704 22836 11756
rect 22888 11744 22894 11756
rect 23474 11744 23480 11756
rect 22888 11716 23480 11744
rect 22888 11704 22894 11716
rect 23474 11704 23480 11716
rect 23532 11744 23538 11756
rect 23845 11747 23903 11753
rect 23845 11744 23857 11747
rect 23532 11716 23857 11744
rect 23532 11704 23538 11716
rect 23845 11713 23857 11716
rect 23891 11713 23903 11747
rect 23845 11707 23903 11713
rect 25774 11704 25780 11756
rect 25832 11704 25838 11756
rect 26326 11704 26332 11756
rect 26384 11704 26390 11756
rect 26421 11747 26479 11753
rect 26421 11713 26433 11747
rect 26467 11713 26479 11747
rect 26421 11707 26479 11713
rect 15105 11679 15163 11685
rect 15105 11676 15117 11679
rect 14056 11648 15117 11676
rect 14056 11636 14062 11648
rect 15105 11645 15117 11648
rect 15151 11645 15163 11679
rect 15105 11639 15163 11645
rect 17681 11679 17739 11685
rect 17681 11645 17693 11679
rect 17727 11645 17739 11679
rect 19153 11679 19211 11685
rect 19153 11676 19165 11679
rect 17681 11639 17739 11645
rect 18984 11648 19165 11676
rect 3712 11580 4384 11608
rect 5445 11543 5503 11549
rect 5445 11509 5457 11543
rect 5491 11540 5503 11543
rect 6730 11540 6736 11552
rect 5491 11512 6736 11540
rect 5491 11509 5503 11512
rect 5445 11503 5503 11509
rect 6730 11500 6736 11512
rect 6788 11500 6794 11552
rect 8389 11543 8447 11549
rect 8389 11509 8401 11543
rect 8435 11540 8447 11543
rect 13078 11540 13084 11552
rect 8435 11512 13084 11540
rect 8435 11509 8447 11512
rect 8389 11503 8447 11509
rect 13078 11500 13084 11512
rect 13136 11500 13142 11552
rect 13909 11543 13967 11549
rect 13909 11509 13921 11543
rect 13955 11540 13967 11543
rect 14090 11540 14096 11552
rect 13955 11512 14096 11540
rect 13955 11509 13967 11512
rect 13909 11503 13967 11509
rect 14090 11500 14096 11512
rect 14148 11500 14154 11552
rect 17696 11540 17724 11639
rect 18984 11552 19012 11648
rect 19153 11645 19165 11648
rect 19199 11645 19211 11679
rect 26436 11676 26464 11707
rect 26694 11704 26700 11756
rect 26752 11744 26758 11756
rect 27525 11747 27583 11753
rect 27525 11744 27537 11747
rect 26752 11716 27537 11744
rect 26752 11704 26758 11716
rect 27525 11713 27537 11716
rect 27571 11713 27583 11747
rect 27525 11707 27583 11713
rect 28074 11676 28080 11688
rect 26436 11648 28080 11676
rect 19153 11639 19211 11645
rect 28074 11636 28080 11648
rect 28132 11636 28138 11688
rect 18966 11540 18972 11552
rect 17696 11512 18972 11540
rect 18966 11500 18972 11512
rect 19024 11500 19030 11552
rect 19061 11543 19119 11549
rect 19061 11509 19073 11543
rect 19107 11540 19119 11543
rect 20346 11540 20352 11552
rect 19107 11512 20352 11540
rect 19107 11509 19119 11512
rect 19061 11503 19119 11509
rect 20346 11500 20352 11512
rect 20404 11500 20410 11552
rect 20533 11543 20591 11549
rect 20533 11509 20545 11543
rect 20579 11540 20591 11543
rect 21082 11540 21088 11552
rect 20579 11512 21088 11540
rect 20579 11509 20591 11512
rect 20533 11503 20591 11509
rect 21082 11500 21088 11512
rect 21140 11500 21146 11552
rect 21174 11500 21180 11552
rect 21232 11540 21238 11552
rect 23382 11540 23388 11552
rect 21232 11512 23388 11540
rect 21232 11500 21238 11512
rect 23382 11500 23388 11512
rect 23440 11500 23446 11552
rect 25590 11500 25596 11552
rect 25648 11500 25654 11552
rect 26145 11543 26203 11549
rect 26145 11509 26157 11543
rect 26191 11540 26203 11543
rect 26418 11540 26424 11552
rect 26191 11512 26424 11540
rect 26191 11509 26203 11512
rect 26145 11503 26203 11509
rect 26418 11500 26424 11512
rect 26476 11500 26482 11552
rect 26510 11500 26516 11552
rect 26568 11540 26574 11552
rect 26973 11543 27031 11549
rect 26973 11540 26985 11543
rect 26568 11512 26985 11540
rect 26568 11500 26574 11512
rect 26973 11509 26985 11512
rect 27019 11509 27031 11543
rect 26973 11503 27031 11509
rect 1104 11450 31832 11472
rect 1104 11398 4182 11450
rect 4234 11398 4246 11450
rect 4298 11398 4310 11450
rect 4362 11398 4374 11450
rect 4426 11398 4438 11450
rect 4490 11398 4502 11450
rect 4554 11398 10182 11450
rect 10234 11398 10246 11450
rect 10298 11398 10310 11450
rect 10362 11398 10374 11450
rect 10426 11398 10438 11450
rect 10490 11398 10502 11450
rect 10554 11398 16182 11450
rect 16234 11398 16246 11450
rect 16298 11398 16310 11450
rect 16362 11398 16374 11450
rect 16426 11398 16438 11450
rect 16490 11398 16502 11450
rect 16554 11398 22182 11450
rect 22234 11398 22246 11450
rect 22298 11398 22310 11450
rect 22362 11398 22374 11450
rect 22426 11398 22438 11450
rect 22490 11398 22502 11450
rect 22554 11398 28182 11450
rect 28234 11398 28246 11450
rect 28298 11398 28310 11450
rect 28362 11398 28374 11450
rect 28426 11398 28438 11450
rect 28490 11398 28502 11450
rect 28554 11398 31832 11450
rect 1104 11376 31832 11398
rect 2590 11336 2596 11348
rect 2240 11308 2596 11336
rect 2133 11271 2191 11277
rect 2133 11237 2145 11271
rect 2179 11237 2191 11271
rect 2133 11231 2191 11237
rect 1949 11135 2007 11141
rect 1949 11101 1961 11135
rect 1995 11101 2007 11135
rect 2148 11132 2176 11231
rect 2240 11209 2268 11308
rect 2590 11296 2596 11308
rect 2648 11296 2654 11348
rect 3694 11296 3700 11348
rect 3752 11336 3758 11348
rect 5537 11339 5595 11345
rect 3752 11308 4292 11336
rect 3752 11296 3758 11308
rect 3789 11271 3847 11277
rect 3789 11237 3801 11271
rect 3835 11237 3847 11271
rect 3789 11231 3847 11237
rect 4264 11268 4292 11308
rect 5537 11305 5549 11339
rect 5583 11336 5595 11339
rect 5626 11336 5632 11348
rect 5583 11308 5632 11336
rect 5583 11305 5595 11308
rect 5537 11299 5595 11305
rect 5626 11296 5632 11308
rect 5684 11296 5690 11348
rect 6178 11296 6184 11348
rect 6236 11336 6242 11348
rect 7374 11336 7380 11348
rect 6236 11308 7380 11336
rect 6236 11296 6242 11308
rect 7374 11296 7380 11308
rect 7432 11296 7438 11348
rect 14090 11296 14096 11348
rect 14148 11296 14154 11348
rect 16022 11296 16028 11348
rect 16080 11296 16086 11348
rect 17954 11296 17960 11348
rect 18012 11336 18018 11348
rect 18049 11339 18107 11345
rect 18049 11336 18061 11339
rect 18012 11308 18061 11336
rect 18012 11296 18018 11308
rect 18049 11305 18061 11308
rect 18095 11305 18107 11339
rect 18049 11299 18107 11305
rect 18785 11339 18843 11345
rect 18785 11305 18797 11339
rect 18831 11336 18843 11339
rect 19426 11336 19432 11348
rect 18831 11308 19432 11336
rect 18831 11305 18843 11308
rect 18785 11299 18843 11305
rect 19426 11296 19432 11308
rect 19484 11296 19490 11348
rect 21266 11296 21272 11348
rect 21324 11336 21330 11348
rect 21913 11339 21971 11345
rect 21913 11336 21925 11339
rect 21324 11308 21925 11336
rect 21324 11296 21330 11308
rect 21913 11305 21925 11308
rect 21959 11305 21971 11339
rect 21913 11299 21971 11305
rect 22741 11339 22799 11345
rect 22741 11305 22753 11339
rect 22787 11336 22799 11339
rect 22830 11336 22836 11348
rect 22787 11308 22836 11336
rect 22787 11305 22799 11308
rect 22741 11299 22799 11305
rect 22830 11296 22836 11308
rect 22888 11296 22894 11348
rect 25222 11296 25228 11348
rect 25280 11296 25286 11348
rect 26605 11339 26663 11345
rect 26605 11305 26617 11339
rect 26651 11336 26663 11339
rect 26694 11336 26700 11348
rect 26651 11308 26700 11336
rect 26651 11305 26663 11308
rect 26605 11299 26663 11305
rect 26694 11296 26700 11308
rect 26752 11296 26758 11348
rect 28074 11296 28080 11348
rect 28132 11296 28138 11348
rect 4264 11240 4752 11268
rect 2225 11203 2283 11209
rect 2225 11169 2237 11203
rect 2271 11169 2283 11203
rect 2225 11163 2283 11169
rect 2481 11135 2539 11141
rect 2481 11132 2493 11135
rect 2148 11104 2493 11132
rect 1949 11095 2007 11101
rect 2481 11101 2493 11104
rect 2527 11101 2539 11135
rect 2481 11095 2539 11101
rect 1964 11064 1992 11095
rect 3804 11064 3832 11231
rect 4062 11160 4068 11212
rect 4120 11160 4126 11212
rect 4264 11209 4292 11240
rect 4249 11203 4307 11209
rect 4249 11169 4261 11203
rect 4295 11169 4307 11203
rect 4249 11163 4307 11169
rect 4341 11203 4399 11209
rect 4341 11169 4353 11203
rect 4387 11169 4399 11203
rect 4724 11200 4752 11240
rect 8570 11228 8576 11280
rect 8628 11268 8634 11280
rect 8757 11271 8815 11277
rect 8757 11268 8769 11271
rect 8628 11240 8769 11268
rect 8628 11228 8634 11240
rect 8757 11237 8769 11240
rect 8803 11268 8815 11271
rect 8803 11240 10548 11268
rect 8803 11237 8815 11240
rect 8757 11231 8815 11237
rect 5902 11200 5908 11212
rect 4724 11172 5908 11200
rect 4341 11163 4399 11169
rect 4080 11132 4108 11160
rect 4356 11132 4384 11163
rect 5902 11160 5908 11172
rect 5960 11160 5966 11212
rect 10520 11209 10548 11240
rect 7377 11203 7435 11209
rect 7377 11200 7389 11203
rect 6932 11172 7389 11200
rect 5166 11132 5172 11144
rect 4080 11104 4384 11132
rect 4724 11104 5172 11132
rect 1964 11036 3832 11064
rect 4157 11067 4215 11073
rect 4157 11033 4169 11067
rect 4203 11064 4215 11067
rect 4617 11067 4675 11073
rect 4617 11064 4629 11067
rect 4203 11036 4629 11064
rect 4203 11033 4215 11036
rect 4157 11027 4215 11033
rect 4617 11033 4629 11036
rect 4663 11033 4675 11067
rect 4617 11027 4675 11033
rect 3605 10999 3663 11005
rect 3605 10965 3617 10999
rect 3651 10996 3663 10999
rect 4724 10996 4752 11104
rect 5166 11092 5172 11104
rect 5224 11092 5230 11144
rect 6362 11092 6368 11144
rect 6420 11132 6426 11144
rect 6932 11141 6960 11172
rect 7377 11169 7389 11172
rect 7423 11169 7435 11203
rect 7377 11163 7435 11169
rect 10505 11203 10563 11209
rect 10505 11169 10517 11203
rect 10551 11169 10563 11203
rect 10505 11163 10563 11169
rect 6917 11135 6975 11141
rect 6917 11132 6929 11135
rect 6420 11104 6929 11132
rect 6420 11092 6426 11104
rect 6917 11101 6929 11104
rect 6963 11101 6975 11135
rect 6917 11095 6975 11101
rect 7098 11092 7104 11144
rect 7156 11132 7162 11144
rect 7193 11135 7251 11141
rect 7193 11132 7205 11135
rect 7156 11104 7205 11132
rect 7156 11092 7162 11104
rect 7193 11101 7205 11104
rect 7239 11101 7251 11135
rect 7392 11132 7420 11163
rect 11330 11160 11336 11212
rect 11388 11200 11394 11212
rect 11701 11203 11759 11209
rect 11701 11200 11713 11203
rect 11388 11172 11713 11200
rect 11388 11160 11394 11172
rect 11701 11169 11713 11172
rect 11747 11169 11759 11203
rect 11701 11163 11759 11169
rect 13722 11160 13728 11212
rect 13780 11200 13786 11212
rect 14108 11200 14136 11296
rect 16040 11200 16068 11296
rect 16114 11228 16120 11280
rect 16172 11268 16178 11280
rect 16301 11271 16359 11277
rect 16301 11268 16313 11271
rect 16172 11240 16313 11268
rect 16172 11228 16178 11240
rect 16301 11237 16313 11240
rect 16347 11237 16359 11271
rect 16301 11231 16359 11237
rect 19245 11271 19303 11277
rect 19245 11237 19257 11271
rect 19291 11237 19303 11271
rect 19245 11231 19303 11237
rect 19904 11240 22600 11268
rect 19260 11200 19288 11231
rect 19904 11209 19932 11240
rect 13780 11172 14044 11200
rect 14108 11172 14228 11200
rect 16040 11172 16528 11200
rect 13780 11160 13786 11172
rect 9030 11132 9036 11144
rect 7392 11104 9036 11132
rect 7193 11095 7251 11101
rect 9030 11092 9036 11104
rect 9088 11092 9094 11144
rect 10873 11135 10931 11141
rect 10873 11101 10885 11135
rect 10919 11132 10931 11135
rect 11514 11132 11520 11144
rect 10919 11104 11520 11132
rect 10919 11101 10931 11104
rect 10873 11095 10931 11101
rect 11514 11092 11520 11104
rect 11572 11092 11578 11144
rect 12986 11132 12992 11144
rect 12406 11104 12992 11132
rect 6672 11067 6730 11073
rect 6672 11033 6684 11067
rect 6718 11064 6730 11067
rect 7644 11067 7702 11073
rect 6718 11036 7052 11064
rect 6718 11033 6730 11036
rect 6672 11027 6730 11033
rect 7024 11005 7052 11036
rect 7644 11033 7656 11067
rect 7690 11064 7702 11067
rect 8478 11064 8484 11076
rect 7690 11036 8484 11064
rect 7690 11033 7702 11036
rect 7644 11027 7702 11033
rect 8478 11024 8484 11036
rect 8536 11024 8542 11076
rect 9858 11024 9864 11076
rect 9916 11064 9922 11076
rect 12406 11064 12434 11104
rect 12986 11092 12992 11104
rect 13044 11132 13050 11144
rect 14016 11132 14044 11172
rect 14090 11132 14096 11144
rect 13044 11104 13860 11132
rect 14016 11104 14096 11132
rect 13044 11092 13050 11104
rect 9916 11036 12434 11064
rect 9916 11024 9922 11036
rect 13722 11024 13728 11076
rect 13780 11024 13786 11076
rect 13832 11008 13860 11104
rect 14090 11092 14096 11104
rect 14148 11092 14154 11144
rect 14200 11132 14228 11172
rect 16500 11141 16528 11172
rect 18248 11172 19288 11200
rect 19889 11203 19947 11209
rect 18248 11141 18276 11172
rect 19889 11169 19901 11203
rect 19935 11169 19947 11203
rect 19889 11163 19947 11169
rect 20346 11160 20352 11212
rect 20404 11200 20410 11212
rect 20717 11203 20775 11209
rect 20717 11200 20729 11203
rect 20404 11172 20729 11200
rect 20404 11160 20410 11172
rect 20717 11169 20729 11172
rect 20763 11200 20775 11203
rect 20763 11172 21404 11200
rect 20763 11169 20775 11172
rect 20717 11163 20775 11169
rect 14349 11135 14407 11141
rect 14349 11132 14361 11135
rect 14200 11104 14361 11132
rect 14349 11101 14361 11104
rect 14395 11101 14407 11135
rect 16117 11135 16175 11141
rect 16117 11132 16129 11135
rect 14349 11095 14407 11101
rect 15488 11104 16129 11132
rect 15488 11008 15516 11104
rect 16117 11101 16129 11104
rect 16163 11101 16175 11135
rect 16117 11095 16175 11101
rect 16485 11135 16543 11141
rect 16485 11101 16497 11135
rect 16531 11101 16543 11135
rect 16485 11095 16543 11101
rect 18233 11135 18291 11141
rect 18233 11101 18245 11135
rect 18279 11101 18291 11135
rect 18233 11095 18291 11101
rect 18601 11135 18659 11141
rect 18601 11101 18613 11135
rect 18647 11132 18659 11135
rect 19242 11132 19248 11144
rect 18647 11104 19248 11132
rect 18647 11101 18659 11104
rect 18601 11095 18659 11101
rect 19242 11092 19248 11104
rect 19300 11092 19306 11144
rect 21376 11141 21404 11172
rect 22094 11160 22100 11212
rect 22152 11160 22158 11212
rect 22572 11209 22600 11240
rect 22557 11203 22615 11209
rect 22557 11169 22569 11203
rect 22603 11200 22615 11203
rect 25240 11200 25268 11296
rect 22603 11172 25268 11200
rect 28092 11200 28120 11296
rect 28721 11203 28779 11209
rect 28721 11200 28733 11203
rect 28092 11172 28733 11200
rect 22603 11169 22615 11172
rect 22557 11163 22615 11169
rect 28721 11169 28733 11172
rect 28767 11169 28779 11203
rect 28721 11163 28779 11169
rect 20993 11135 21051 11141
rect 20993 11101 21005 11135
rect 21039 11132 21051 11135
rect 21361 11135 21419 11141
rect 21039 11104 21312 11132
rect 21039 11101 21051 11104
rect 20993 11095 21051 11101
rect 19613 11067 19671 11073
rect 19613 11033 19625 11067
rect 19659 11064 19671 11067
rect 20073 11067 20131 11073
rect 20073 11064 20085 11067
rect 19659 11036 20085 11064
rect 19659 11033 19671 11036
rect 19613 11027 19671 11033
rect 20073 11033 20085 11036
rect 20119 11033 20131 11067
rect 20073 11027 20131 11033
rect 21082 11024 21088 11076
rect 21140 11024 21146 11076
rect 21174 11024 21180 11076
rect 21232 11024 21238 11076
rect 21284 11064 21312 11104
rect 21361 11101 21373 11135
rect 21407 11101 21419 11135
rect 22112 11132 22140 11160
rect 22281 11135 22339 11141
rect 22281 11132 22293 11135
rect 22112 11104 22293 11132
rect 21361 11095 21419 11101
rect 22281 11101 22293 11104
rect 22327 11101 22339 11135
rect 22281 11095 22339 11101
rect 22738 11092 22744 11144
rect 22796 11132 22802 11144
rect 22925 11135 22983 11141
rect 22925 11132 22937 11135
rect 22796 11104 22937 11132
rect 22796 11092 22802 11104
rect 22925 11101 22937 11104
rect 22971 11101 22983 11135
rect 22925 11095 22983 11101
rect 23017 11135 23075 11141
rect 23017 11101 23029 11135
rect 23063 11132 23075 11135
rect 23293 11135 23351 11141
rect 23063 11104 23244 11132
rect 23063 11101 23075 11104
rect 23017 11095 23075 11101
rect 22756 11064 22784 11092
rect 21284 11036 22784 11064
rect 23106 11024 23112 11076
rect 23164 11024 23170 11076
rect 23216 11064 23244 11104
rect 23293 11101 23305 11135
rect 23339 11132 23351 11135
rect 23474 11132 23480 11144
rect 23339 11104 23480 11132
rect 23339 11101 23351 11104
rect 23293 11095 23351 11101
rect 23474 11092 23480 11104
rect 23532 11092 23538 11144
rect 23842 11092 23848 11144
rect 23900 11092 23906 11144
rect 25222 11092 25228 11144
rect 25280 11132 25286 11144
rect 26050 11132 26056 11144
rect 25280 11104 26056 11132
rect 25280 11092 25286 11104
rect 26050 11092 26056 11104
rect 26108 11132 26114 11144
rect 26697 11135 26755 11141
rect 26697 11132 26709 11135
rect 26108 11104 26709 11132
rect 26108 11092 26114 11104
rect 26697 11101 26709 11104
rect 26743 11101 26755 11135
rect 26697 11095 26755 11101
rect 23860 11064 23888 11092
rect 23216 11036 23888 11064
rect 25492 11067 25550 11073
rect 25492 11033 25504 11067
rect 25538 11064 25550 11067
rect 25590 11064 25596 11076
rect 25538 11036 25596 11064
rect 25538 11033 25550 11036
rect 25492 11027 25550 11033
rect 25590 11024 25596 11036
rect 25648 11024 25654 11076
rect 26786 11024 26792 11076
rect 26844 11064 26850 11076
rect 26942 11067 27000 11073
rect 26942 11064 26954 11067
rect 26844 11036 26954 11064
rect 26844 11024 26850 11036
rect 26942 11033 26954 11036
rect 26988 11033 27000 11067
rect 26942 11027 27000 11033
rect 3651 10968 4752 10996
rect 7009 10999 7067 11005
rect 3651 10965 3663 10968
rect 3605 10959 3663 10965
rect 7009 10965 7021 10999
rect 7055 10965 7067 10999
rect 7009 10959 7067 10965
rect 9950 10956 9956 11008
rect 10008 10956 10014 11008
rect 10686 10956 10692 11008
rect 10744 10956 10750 11008
rect 12342 10956 12348 11008
rect 12400 10956 12406 11008
rect 13814 10956 13820 11008
rect 13872 10956 13878 11008
rect 15470 10956 15476 11008
rect 15528 10956 15534 11008
rect 15562 10956 15568 11008
rect 15620 10956 15626 11008
rect 19426 10956 19432 11008
rect 19484 10996 19490 11008
rect 19702 10996 19708 11008
rect 19484 10968 19708 10996
rect 19484 10956 19490 10968
rect 19702 10956 19708 10968
rect 19760 10956 19766 11008
rect 20806 10956 20812 11008
rect 20864 10956 20870 11008
rect 22373 10999 22431 11005
rect 22373 10965 22385 10999
rect 22419 10996 22431 10999
rect 24670 10996 24676 11008
rect 22419 10968 24676 10996
rect 22419 10965 22431 10968
rect 22373 10959 22431 10965
rect 24670 10956 24676 10968
rect 24728 10956 24734 11008
rect 28166 10956 28172 11008
rect 28224 10956 28230 11008
rect 1104 10906 31832 10928
rect 1104 10854 4922 10906
rect 4974 10854 4986 10906
rect 5038 10854 5050 10906
rect 5102 10854 5114 10906
rect 5166 10854 5178 10906
rect 5230 10854 5242 10906
rect 5294 10854 10922 10906
rect 10974 10854 10986 10906
rect 11038 10854 11050 10906
rect 11102 10854 11114 10906
rect 11166 10854 11178 10906
rect 11230 10854 11242 10906
rect 11294 10854 16922 10906
rect 16974 10854 16986 10906
rect 17038 10854 17050 10906
rect 17102 10854 17114 10906
rect 17166 10854 17178 10906
rect 17230 10854 17242 10906
rect 17294 10854 22922 10906
rect 22974 10854 22986 10906
rect 23038 10854 23050 10906
rect 23102 10854 23114 10906
rect 23166 10854 23178 10906
rect 23230 10854 23242 10906
rect 23294 10854 28922 10906
rect 28974 10854 28986 10906
rect 29038 10854 29050 10906
rect 29102 10854 29114 10906
rect 29166 10854 29178 10906
rect 29230 10854 29242 10906
rect 29294 10854 31832 10906
rect 1104 10832 31832 10854
rect 6089 10795 6147 10801
rect 6089 10761 6101 10795
rect 6135 10761 6147 10795
rect 6089 10755 6147 10761
rect 4433 10727 4491 10733
rect 4433 10693 4445 10727
rect 4479 10724 4491 10727
rect 4706 10724 4712 10736
rect 4479 10696 4712 10724
rect 4479 10693 4491 10696
rect 4433 10687 4491 10693
rect 4706 10684 4712 10696
rect 4764 10684 4770 10736
rect 5813 10727 5871 10733
rect 5813 10724 5825 10727
rect 5184 10696 5825 10724
rect 5184 10668 5212 10696
rect 5813 10693 5825 10696
rect 5859 10693 5871 10727
rect 5813 10687 5871 10693
rect 2590 10616 2596 10668
rect 2648 10656 2654 10668
rect 2757 10659 2815 10665
rect 2757 10656 2769 10659
rect 2648 10628 2769 10656
rect 2648 10616 2654 10628
rect 2757 10625 2769 10628
rect 2803 10625 2815 10659
rect 2757 10619 2815 10625
rect 4341 10659 4399 10665
rect 4341 10625 4353 10659
rect 4387 10656 4399 10659
rect 4801 10659 4859 10665
rect 4801 10656 4813 10659
rect 4387 10628 4813 10656
rect 4387 10625 4399 10628
rect 4341 10619 4399 10625
rect 4801 10625 4813 10628
rect 4847 10625 4859 10659
rect 4801 10619 4859 10625
rect 5166 10616 5172 10668
rect 5224 10616 5230 10668
rect 5537 10659 5595 10665
rect 5537 10625 5549 10659
rect 5583 10625 5595 10659
rect 5537 10619 5595 10625
rect 2498 10548 2504 10600
rect 2556 10548 2562 10600
rect 4614 10548 4620 10600
rect 4672 10548 4678 10600
rect 5353 10591 5411 10597
rect 5353 10557 5365 10591
rect 5399 10588 5411 10591
rect 5552 10588 5580 10619
rect 5626 10616 5632 10668
rect 5684 10656 5690 10668
rect 5721 10659 5779 10665
rect 5721 10656 5733 10659
rect 5684 10628 5733 10656
rect 5684 10616 5690 10628
rect 5721 10625 5733 10628
rect 5767 10625 5779 10659
rect 5721 10619 5779 10625
rect 5905 10659 5963 10665
rect 5905 10625 5917 10659
rect 5951 10625 5963 10659
rect 6104 10656 6132 10755
rect 6914 10752 6920 10804
rect 6972 10752 6978 10804
rect 7006 10752 7012 10804
rect 7064 10792 7070 10804
rect 7285 10795 7343 10801
rect 7285 10792 7297 10795
rect 7064 10764 7297 10792
rect 7064 10752 7070 10764
rect 7285 10761 7297 10764
rect 7331 10761 7343 10795
rect 7285 10755 7343 10761
rect 8205 10795 8263 10801
rect 8205 10761 8217 10795
rect 8251 10792 8263 10795
rect 8386 10792 8392 10804
rect 8251 10764 8392 10792
rect 8251 10761 8263 10764
rect 8205 10755 8263 10761
rect 8386 10752 8392 10764
rect 8444 10752 8450 10804
rect 8481 10795 8539 10801
rect 8481 10761 8493 10795
rect 8527 10792 8539 10795
rect 8570 10792 8576 10804
rect 8527 10764 8576 10792
rect 8527 10761 8539 10764
rect 8481 10755 8539 10761
rect 8570 10752 8576 10764
rect 8628 10752 8634 10804
rect 8662 10752 8668 10804
rect 8720 10792 8726 10804
rect 8941 10795 8999 10801
rect 8941 10792 8953 10795
rect 8720 10764 8953 10792
rect 8720 10752 8726 10764
rect 8941 10761 8953 10764
rect 8987 10761 8999 10795
rect 8941 10755 8999 10761
rect 9309 10795 9367 10801
rect 9309 10761 9321 10795
rect 9355 10792 9367 10795
rect 9950 10792 9956 10804
rect 9355 10764 9956 10792
rect 9355 10761 9367 10764
rect 9309 10755 9367 10761
rect 9950 10752 9956 10764
rect 10008 10752 10014 10804
rect 11330 10752 11336 10804
rect 11388 10752 11394 10804
rect 11514 10752 11520 10804
rect 11572 10752 11578 10804
rect 11885 10795 11943 10801
rect 11885 10761 11897 10795
rect 11931 10792 11943 10795
rect 12342 10792 12348 10804
rect 11931 10764 12348 10792
rect 11931 10761 11943 10764
rect 11885 10755 11943 10761
rect 12342 10752 12348 10764
rect 12400 10752 12406 10804
rect 14182 10752 14188 10804
rect 14240 10752 14246 10804
rect 14553 10795 14611 10801
rect 14553 10761 14565 10795
rect 14599 10792 14611 10795
rect 15562 10792 15568 10804
rect 14599 10764 15568 10792
rect 14599 10761 14611 10764
rect 14553 10755 14611 10761
rect 15562 10752 15568 10764
rect 15620 10752 15626 10804
rect 25685 10795 25743 10801
rect 25685 10761 25697 10795
rect 25731 10792 25743 10795
rect 25774 10792 25780 10804
rect 25731 10764 25780 10792
rect 25731 10761 25743 10764
rect 25685 10755 25743 10761
rect 25774 10752 25780 10764
rect 25832 10752 25838 10804
rect 26053 10795 26111 10801
rect 26053 10761 26065 10795
rect 26099 10792 26111 10795
rect 26510 10792 26516 10804
rect 26099 10764 26516 10792
rect 26099 10761 26111 10764
rect 26053 10755 26111 10761
rect 26510 10752 26516 10764
rect 26568 10752 26574 10804
rect 26697 10795 26755 10801
rect 26697 10761 26709 10795
rect 26743 10792 26755 10795
rect 26786 10792 26792 10804
rect 26743 10764 26792 10792
rect 26743 10761 26755 10764
rect 26697 10755 26755 10761
rect 26786 10752 26792 10764
rect 26844 10752 26850 10804
rect 27341 10795 27399 10801
rect 27341 10761 27353 10795
rect 27387 10792 27399 10795
rect 28166 10792 28172 10804
rect 27387 10764 28172 10792
rect 27387 10761 27399 10764
rect 27341 10755 27399 10761
rect 28166 10752 28172 10764
rect 28224 10752 28230 10804
rect 29362 10792 29368 10804
rect 28966 10764 29368 10792
rect 6825 10727 6883 10733
rect 6825 10693 6837 10727
rect 6871 10724 6883 10727
rect 7190 10724 7196 10736
rect 6871 10696 7196 10724
rect 6871 10693 6883 10696
rect 6825 10687 6883 10693
rect 7190 10684 7196 10696
rect 7248 10684 7254 10736
rect 10220 10727 10278 10733
rect 8220 10696 8524 10724
rect 8021 10659 8079 10665
rect 8021 10656 8033 10659
rect 6104 10628 8033 10656
rect 5905 10619 5963 10625
rect 8021 10625 8033 10628
rect 8067 10625 8079 10659
rect 8021 10619 8079 10625
rect 5399 10560 5580 10588
rect 5920 10588 5948 10619
rect 6178 10588 6184 10600
rect 5920 10560 6184 10588
rect 5399 10557 5411 10560
rect 5353 10551 5411 10557
rect 3881 10523 3939 10529
rect 3881 10489 3893 10523
rect 3927 10520 3939 10523
rect 5368 10520 5396 10551
rect 6178 10548 6184 10560
rect 6236 10548 6242 10600
rect 6641 10591 6699 10597
rect 6641 10588 6653 10591
rect 6288 10560 6653 10588
rect 3927 10492 5396 10520
rect 3927 10489 3939 10492
rect 3881 10483 3939 10489
rect 3970 10412 3976 10464
rect 4028 10412 4034 10464
rect 4062 10412 4068 10464
rect 4120 10452 4126 10464
rect 6288 10452 6316 10560
rect 6641 10557 6653 10560
rect 6687 10557 6699 10591
rect 6641 10551 6699 10557
rect 6730 10548 6736 10600
rect 6788 10588 6794 10600
rect 8220 10588 8248 10696
rect 8297 10659 8355 10665
rect 8297 10625 8309 10659
rect 8343 10656 8355 10659
rect 8389 10659 8447 10665
rect 8389 10656 8401 10659
rect 8343 10628 8401 10656
rect 8343 10625 8355 10628
rect 8297 10619 8355 10625
rect 8389 10625 8401 10628
rect 8435 10625 8447 10659
rect 8496 10656 8524 10696
rect 10220 10693 10232 10727
rect 10266 10724 10278 10727
rect 10686 10724 10692 10736
rect 10266 10696 10692 10724
rect 10266 10693 10278 10696
rect 10220 10687 10278 10693
rect 10686 10684 10692 10696
rect 10744 10684 10750 10736
rect 10870 10684 10876 10736
rect 10928 10684 10934 10736
rect 11606 10684 11612 10736
rect 11664 10724 11670 10736
rect 12989 10727 13047 10733
rect 12989 10724 13001 10727
rect 11664 10696 13001 10724
rect 11664 10684 11670 10696
rect 12989 10693 13001 10696
rect 13035 10693 13047 10727
rect 12989 10687 13047 10693
rect 13814 10684 13820 10736
rect 13872 10684 13878 10736
rect 24394 10684 24400 10736
rect 24452 10724 24458 10736
rect 28966 10724 28994 10764
rect 29362 10752 29368 10764
rect 29420 10792 29426 10804
rect 29730 10792 29736 10804
rect 29420 10764 29736 10792
rect 29420 10752 29426 10764
rect 29730 10752 29736 10764
rect 29788 10752 29794 10804
rect 24452 10696 28994 10724
rect 24452 10684 24458 10696
rect 8665 10659 8723 10665
rect 8665 10656 8677 10659
rect 8496 10628 8677 10656
rect 8389 10619 8447 10625
rect 8665 10625 8677 10628
rect 8711 10625 8723 10659
rect 8665 10619 8723 10625
rect 9401 10659 9459 10665
rect 9401 10625 9413 10659
rect 9447 10656 9459 10659
rect 10888 10656 10916 10684
rect 11977 10659 12035 10665
rect 11977 10656 11989 10659
rect 9447 10628 11989 10656
rect 9447 10625 9459 10628
rect 9401 10619 9459 10625
rect 11977 10625 11989 10628
rect 12023 10625 12035 10659
rect 11977 10619 12035 10625
rect 14645 10659 14703 10665
rect 14645 10625 14657 10659
rect 14691 10656 14703 10659
rect 15102 10656 15108 10668
rect 14691 10628 15108 10656
rect 14691 10625 14703 10628
rect 14645 10619 14703 10625
rect 6788 10560 8248 10588
rect 8404 10588 8432 10619
rect 15102 10616 15108 10628
rect 15160 10616 15166 10668
rect 19518 10616 19524 10668
rect 19576 10656 19582 10668
rect 19613 10659 19671 10665
rect 19613 10656 19625 10659
rect 19576 10628 19625 10656
rect 19576 10616 19582 10628
rect 19613 10625 19625 10628
rect 19659 10625 19671 10659
rect 19613 10619 19671 10625
rect 19889 10659 19947 10665
rect 19889 10625 19901 10659
rect 19935 10656 19947 10659
rect 20254 10656 20260 10668
rect 19935 10628 20260 10656
rect 19935 10625 19947 10628
rect 19889 10619 19947 10625
rect 20254 10616 20260 10628
rect 20312 10616 20318 10668
rect 20346 10616 20352 10668
rect 20404 10616 20410 10668
rect 26513 10659 26571 10665
rect 25332 10628 26280 10656
rect 25332 10600 25360 10628
rect 8404 10560 8524 10588
rect 6788 10548 6794 10560
rect 8496 10520 8524 10560
rect 8570 10548 8576 10600
rect 8628 10588 8634 10600
rect 9493 10591 9551 10597
rect 9493 10588 9505 10591
rect 8628 10560 9505 10588
rect 8628 10548 8634 10560
rect 9493 10557 9505 10560
rect 9539 10557 9551 10591
rect 9493 10551 9551 10557
rect 9953 10591 10011 10597
rect 9953 10557 9965 10591
rect 9999 10557 10011 10591
rect 9953 10551 10011 10557
rect 8496 10492 8984 10520
rect 4120 10424 6316 10452
rect 7837 10455 7895 10461
rect 4120 10412 4126 10424
rect 7837 10421 7849 10455
rect 7883 10452 7895 10455
rect 8754 10452 8760 10464
rect 7883 10424 8760 10452
rect 7883 10421 7895 10424
rect 7837 10415 7895 10421
rect 8754 10412 8760 10424
rect 8812 10412 8818 10464
rect 8846 10412 8852 10464
rect 8904 10412 8910 10464
rect 8956 10452 8984 10492
rect 9030 10480 9036 10532
rect 9088 10520 9094 10532
rect 9968 10520 9996 10551
rect 12158 10548 12164 10600
rect 12216 10548 12222 10600
rect 14829 10591 14887 10597
rect 14829 10557 14841 10591
rect 14875 10588 14887 10591
rect 15286 10588 15292 10600
rect 14875 10560 15292 10588
rect 14875 10557 14887 10560
rect 14829 10551 14887 10557
rect 15286 10548 15292 10560
rect 15344 10548 15350 10600
rect 19702 10548 19708 10600
rect 19760 10548 19766 10600
rect 25314 10548 25320 10600
rect 25372 10548 25378 10600
rect 26252 10597 26280 10628
rect 26513 10625 26525 10659
rect 26559 10656 26571 10659
rect 26559 10628 27016 10656
rect 26559 10625 26571 10628
rect 26513 10619 26571 10625
rect 26145 10591 26203 10597
rect 26145 10557 26157 10591
rect 26191 10557 26203 10591
rect 26145 10551 26203 10557
rect 26237 10591 26295 10597
rect 26237 10557 26249 10591
rect 26283 10557 26295 10591
rect 26237 10551 26295 10557
rect 9088 10492 9996 10520
rect 19904 10492 20852 10520
rect 9088 10480 9094 10492
rect 14090 10452 14096 10464
rect 8956 10424 14096 10452
rect 14090 10412 14096 10424
rect 14148 10452 14154 10464
rect 14826 10452 14832 10464
rect 14148 10424 14832 10452
rect 14148 10412 14154 10424
rect 14826 10412 14832 10424
rect 14884 10412 14890 10464
rect 19904 10461 19932 10492
rect 20824 10464 20852 10492
rect 19889 10455 19947 10461
rect 19889 10421 19901 10455
rect 19935 10421 19947 10455
rect 19889 10415 19947 10421
rect 20070 10412 20076 10464
rect 20128 10412 20134 10464
rect 20162 10412 20168 10464
rect 20220 10412 20226 10464
rect 20806 10412 20812 10464
rect 20864 10412 20870 10464
rect 26160 10452 26188 10551
rect 26988 10529 27016 10628
rect 27430 10548 27436 10600
rect 27488 10548 27494 10600
rect 27522 10548 27528 10600
rect 27580 10548 27586 10600
rect 29917 10591 29975 10597
rect 29917 10557 29929 10591
rect 29963 10588 29975 10591
rect 30190 10588 30196 10600
rect 29963 10560 30196 10588
rect 29963 10557 29975 10560
rect 29917 10551 29975 10557
rect 30190 10548 30196 10560
rect 30248 10548 30254 10600
rect 26973 10523 27031 10529
rect 26973 10489 26985 10523
rect 27019 10489 27031 10523
rect 26973 10483 27031 10489
rect 27448 10452 27476 10548
rect 26160 10424 27476 10452
rect 28994 10412 29000 10464
rect 29052 10452 29058 10464
rect 29273 10455 29331 10461
rect 29273 10452 29285 10455
rect 29052 10424 29285 10452
rect 29052 10412 29058 10424
rect 29273 10421 29285 10424
rect 29319 10421 29331 10455
rect 29273 10415 29331 10421
rect 1104 10362 31832 10384
rect 1104 10310 4182 10362
rect 4234 10310 4246 10362
rect 4298 10310 4310 10362
rect 4362 10310 4374 10362
rect 4426 10310 4438 10362
rect 4490 10310 4502 10362
rect 4554 10310 10182 10362
rect 10234 10310 10246 10362
rect 10298 10310 10310 10362
rect 10362 10310 10374 10362
rect 10426 10310 10438 10362
rect 10490 10310 10502 10362
rect 10554 10310 16182 10362
rect 16234 10310 16246 10362
rect 16298 10310 16310 10362
rect 16362 10310 16374 10362
rect 16426 10310 16438 10362
rect 16490 10310 16502 10362
rect 16554 10310 22182 10362
rect 22234 10310 22246 10362
rect 22298 10310 22310 10362
rect 22362 10310 22374 10362
rect 22426 10310 22438 10362
rect 22490 10310 22502 10362
rect 22554 10310 28182 10362
rect 28234 10310 28246 10362
rect 28298 10310 28310 10362
rect 28362 10310 28374 10362
rect 28426 10310 28438 10362
rect 28490 10310 28502 10362
rect 28554 10310 31832 10362
rect 1104 10288 31832 10310
rect 2590 10208 2596 10260
rect 2648 10208 2654 10260
rect 3970 10208 3976 10260
rect 4028 10208 4034 10260
rect 8478 10208 8484 10260
rect 8536 10208 8542 10260
rect 8846 10208 8852 10260
rect 8904 10208 8910 10260
rect 9953 10251 10011 10257
rect 9953 10217 9965 10251
rect 9999 10248 10011 10251
rect 10042 10248 10048 10260
rect 9999 10220 10048 10248
rect 9999 10217 10011 10220
rect 9953 10211 10011 10217
rect 10042 10208 10048 10220
rect 10100 10208 10106 10260
rect 20070 10248 20076 10260
rect 12268 10220 20076 10248
rect 2777 10047 2835 10053
rect 2777 10013 2789 10047
rect 2823 10044 2835 10047
rect 3988 10044 4016 10208
rect 4062 10072 4068 10124
rect 4120 10112 4126 10124
rect 8496 10121 8524 10208
rect 8864 10180 8892 10208
rect 10229 10183 10287 10189
rect 10229 10180 10241 10183
rect 8864 10152 10241 10180
rect 10229 10149 10241 10152
rect 10275 10149 10287 10183
rect 10229 10143 10287 10149
rect 4341 10115 4399 10121
rect 4341 10112 4353 10115
rect 4120 10084 4353 10112
rect 4120 10072 4126 10084
rect 4341 10081 4353 10084
rect 4387 10081 4399 10115
rect 4341 10075 4399 10081
rect 8481 10115 8539 10121
rect 8481 10081 8493 10115
rect 8527 10081 8539 10115
rect 12268 10112 12296 10220
rect 20070 10208 20076 10220
rect 20128 10208 20134 10260
rect 20254 10208 20260 10260
rect 20312 10248 20318 10260
rect 20901 10251 20959 10257
rect 20901 10248 20913 10251
rect 20312 10220 20913 10248
rect 20312 10208 20318 10220
rect 20901 10217 20913 10220
rect 20947 10217 20959 10251
rect 20901 10211 20959 10217
rect 23750 10208 23756 10260
rect 23808 10248 23814 10260
rect 29914 10248 29920 10260
rect 23808 10220 29920 10248
rect 23808 10208 23814 10220
rect 29914 10208 29920 10220
rect 29972 10208 29978 10260
rect 23845 10183 23903 10189
rect 19996 10152 22094 10180
rect 15470 10112 15476 10124
rect 8481 10075 8539 10081
rect 10152 10084 12296 10112
rect 13096 10084 14412 10112
rect 2823 10016 4016 10044
rect 2823 10013 2835 10016
rect 2777 10007 2835 10013
rect 4706 10004 4712 10056
rect 4764 10044 4770 10056
rect 5166 10044 5172 10056
rect 4764 10016 5172 10044
rect 4764 10004 4770 10016
rect 5166 10004 5172 10016
rect 5224 10004 5230 10056
rect 8386 10004 8392 10056
rect 8444 10044 8450 10056
rect 10152 10053 10180 10084
rect 13096 10056 13124 10084
rect 9493 10047 9551 10053
rect 9493 10044 9505 10047
rect 8444 10016 9505 10044
rect 8444 10004 8450 10016
rect 9493 10013 9505 10016
rect 9539 10013 9551 10047
rect 9493 10007 9551 10013
rect 10137 10047 10195 10053
rect 10137 10013 10149 10047
rect 10183 10013 10195 10047
rect 10137 10007 10195 10013
rect 10321 10047 10379 10053
rect 10321 10013 10333 10047
rect 10367 10013 10379 10047
rect 10321 10007 10379 10013
rect 10413 10047 10471 10053
rect 10413 10013 10425 10047
rect 10459 10044 10471 10047
rect 10781 10047 10839 10053
rect 10781 10044 10793 10047
rect 10459 10016 10793 10044
rect 10459 10013 10471 10016
rect 10413 10007 10471 10013
rect 10781 10013 10793 10016
rect 10827 10013 10839 10047
rect 10781 10007 10839 10013
rect 10965 10047 11023 10053
rect 10965 10013 10977 10047
rect 11011 10044 11023 10047
rect 11330 10044 11336 10056
rect 11011 10016 11336 10044
rect 11011 10013 11023 10016
rect 10965 10007 11023 10013
rect 4157 9979 4215 9985
rect 4157 9945 4169 9979
rect 4203 9976 4215 9979
rect 4617 9979 4675 9985
rect 4617 9976 4629 9979
rect 4203 9948 4629 9976
rect 4203 9945 4215 9948
rect 4157 9939 4215 9945
rect 4617 9945 4629 9948
rect 4663 9945 4675 9979
rect 4617 9939 4675 9945
rect 8297 9979 8355 9985
rect 8297 9945 8309 9979
rect 8343 9976 8355 9979
rect 8941 9979 8999 9985
rect 8941 9976 8953 9979
rect 8343 9948 8953 9976
rect 8343 9945 8355 9948
rect 8297 9939 8355 9945
rect 8941 9945 8953 9948
rect 8987 9945 8999 9979
rect 8941 9939 8999 9945
rect 9858 9936 9864 9988
rect 9916 9976 9922 9988
rect 10336 9976 10364 10007
rect 11330 10004 11336 10016
rect 11388 10004 11394 10056
rect 11701 10047 11759 10053
rect 11701 10013 11713 10047
rect 11747 10044 11759 10047
rect 12894 10044 12900 10056
rect 11747 10016 12900 10044
rect 11747 10013 11759 10016
rect 11701 10007 11759 10013
rect 12894 10004 12900 10016
rect 12952 10004 12958 10056
rect 13078 10004 13084 10056
rect 13136 10004 13142 10056
rect 14090 10004 14096 10056
rect 14148 10004 14154 10056
rect 14384 10053 14412 10084
rect 14476 10084 15476 10112
rect 14369 10047 14427 10053
rect 14369 10013 14381 10047
rect 14415 10013 14427 10047
rect 14369 10007 14427 10013
rect 9916 9948 10364 9976
rect 11149 9979 11207 9985
rect 9916 9936 9922 9948
rect 11149 9945 11161 9979
rect 11195 9976 11207 9979
rect 11790 9976 11796 9988
rect 11195 9948 11796 9976
rect 11195 9945 11207 9948
rect 11149 9939 11207 9945
rect 11790 9936 11796 9948
rect 11848 9976 11854 9988
rect 11885 9979 11943 9985
rect 11885 9976 11897 9979
rect 11848 9948 11897 9976
rect 11848 9936 11854 9948
rect 11885 9945 11897 9948
rect 11931 9945 11943 9979
rect 11885 9939 11943 9945
rect 14185 9979 14243 9985
rect 14185 9945 14197 9979
rect 14231 9976 14243 9979
rect 14476 9976 14504 10084
rect 15470 10072 15476 10084
rect 15528 10072 15534 10124
rect 19996 10121 20024 10152
rect 19981 10115 20039 10121
rect 19981 10081 19993 10115
rect 20027 10081 20039 10115
rect 22066 10112 22094 10152
rect 23845 10149 23857 10183
rect 23891 10180 23903 10183
rect 25038 10180 25044 10192
rect 23891 10152 25044 10180
rect 23891 10149 23903 10152
rect 23845 10143 23903 10149
rect 25038 10140 25044 10152
rect 25096 10140 25102 10192
rect 29549 10183 29607 10189
rect 29549 10149 29561 10183
rect 29595 10149 29607 10183
rect 29932 10180 29960 10208
rect 29932 10152 30604 10180
rect 29549 10143 29607 10149
rect 24578 10112 24584 10124
rect 19981 10075 20039 10081
rect 20732 10084 21220 10112
rect 22066 10084 24584 10112
rect 14826 10004 14832 10056
rect 14884 10004 14890 10056
rect 20254 10004 20260 10056
rect 20312 10044 20318 10056
rect 20732 10053 20760 10084
rect 20717 10047 20775 10053
rect 20717 10044 20729 10047
rect 20312 10016 20729 10044
rect 20312 10004 20318 10016
rect 20717 10013 20729 10016
rect 20763 10013 20775 10047
rect 20717 10007 20775 10013
rect 21080 10047 21138 10053
rect 21080 10013 21092 10047
rect 21126 10013 21138 10047
rect 21192 10044 21220 10084
rect 24578 10072 24584 10084
rect 24636 10072 24642 10124
rect 24949 10115 25007 10121
rect 24949 10081 24961 10115
rect 24995 10081 25007 10115
rect 24949 10075 25007 10081
rect 21397 10047 21455 10053
rect 21397 10044 21409 10047
rect 21192 10016 21409 10044
rect 21080 10007 21138 10013
rect 21397 10013 21409 10016
rect 21443 10013 21455 10047
rect 21397 10007 21455 10013
rect 21545 10047 21603 10053
rect 21545 10013 21557 10047
rect 21591 10044 21603 10047
rect 23661 10047 23719 10053
rect 21591 10016 22094 10044
rect 21591 10013 21603 10016
rect 21545 10007 21603 10013
rect 14231 9948 14504 9976
rect 14553 9979 14611 9985
rect 14231 9945 14243 9948
rect 14185 9939 14243 9945
rect 14553 9945 14565 9979
rect 14599 9976 14611 9979
rect 14918 9976 14924 9988
rect 14599 9948 14924 9976
rect 14599 9945 14611 9948
rect 14553 9939 14611 9945
rect 14918 9936 14924 9948
rect 14976 9936 14982 9988
rect 19705 9979 19763 9985
rect 19705 9945 19717 9979
rect 19751 9976 19763 9979
rect 20165 9979 20223 9985
rect 20165 9976 20177 9979
rect 19751 9948 20177 9976
rect 19751 9945 19763 9948
rect 19705 9939 19763 9945
rect 20165 9945 20177 9948
rect 20211 9945 20223 9979
rect 20165 9939 20223 9945
rect 3786 9868 3792 9920
rect 3844 9868 3850 9920
rect 4249 9911 4307 9917
rect 4249 9877 4261 9911
rect 4295 9908 4307 9911
rect 4522 9908 4528 9920
rect 4295 9880 4528 9908
rect 4295 9877 4307 9880
rect 4249 9871 4307 9877
rect 4522 9868 4528 9880
rect 4580 9868 4586 9920
rect 7926 9868 7932 9920
rect 7984 9868 7990 9920
rect 8389 9911 8447 9917
rect 8389 9877 8401 9911
rect 8435 9908 8447 9911
rect 8570 9908 8576 9920
rect 8435 9880 8576 9908
rect 8435 9877 8447 9880
rect 8389 9871 8447 9877
rect 8570 9868 8576 9880
rect 8628 9868 8634 9920
rect 11514 9868 11520 9920
rect 11572 9868 11578 9920
rect 14642 9868 14648 9920
rect 14700 9868 14706 9920
rect 19334 9868 19340 9920
rect 19392 9868 19398 9920
rect 19426 9868 19432 9920
rect 19484 9908 19490 9920
rect 19797 9911 19855 9917
rect 19797 9908 19809 9911
rect 19484 9880 19809 9908
rect 19484 9868 19490 9880
rect 19797 9877 19809 9880
rect 19843 9877 19855 9911
rect 21100 9908 21128 10007
rect 21174 9936 21180 9988
rect 21232 9936 21238 9988
rect 21266 9936 21272 9988
rect 21324 9936 21330 9988
rect 22066 9976 22094 10016
rect 23661 10013 23673 10047
rect 23707 10044 23719 10047
rect 23707 10016 24440 10044
rect 23707 10013 23719 10016
rect 23661 10007 23719 10013
rect 24302 9976 24308 9988
rect 22066 9948 24308 9976
rect 24302 9936 24308 9948
rect 24360 9936 24366 9988
rect 23750 9908 23756 9920
rect 21100 9880 23756 9908
rect 19797 9871 19855 9877
rect 23750 9868 23756 9880
rect 23808 9868 23814 9920
rect 24412 9917 24440 10016
rect 24486 10004 24492 10056
rect 24544 10044 24550 10056
rect 24964 10044 24992 10075
rect 25869 10047 25927 10053
rect 24544 10016 25820 10044
rect 24544 10004 24550 10016
rect 24765 9979 24823 9985
rect 24765 9945 24777 9979
rect 24811 9976 24823 9979
rect 25225 9979 25283 9985
rect 25225 9976 25237 9979
rect 24811 9948 25237 9976
rect 24811 9945 24823 9948
rect 24765 9939 24823 9945
rect 25225 9945 25237 9948
rect 25271 9945 25283 9979
rect 25792 9976 25820 10016
rect 25869 10013 25881 10047
rect 25915 10044 25927 10047
rect 26050 10044 26056 10056
rect 25915 10016 26056 10044
rect 25915 10013 25927 10016
rect 25869 10007 25927 10013
rect 26050 10004 26056 10016
rect 26108 10004 26114 10056
rect 29089 10047 29147 10053
rect 29089 10013 29101 10047
rect 29135 10044 29147 10047
rect 29564 10044 29592 10143
rect 30098 10112 30104 10124
rect 29135 10016 29592 10044
rect 29656 10084 30104 10112
rect 29135 10013 29147 10016
rect 29089 10007 29147 10013
rect 29656 9976 29684 10084
rect 30098 10072 30104 10084
rect 30156 10072 30162 10124
rect 30190 10072 30196 10124
rect 30248 10112 30254 10124
rect 30248 10084 30512 10112
rect 30248 10072 30254 10084
rect 29730 10004 29736 10056
rect 29788 10044 29794 10056
rect 30484 10053 30512 10084
rect 30377 10047 30435 10053
rect 30377 10044 30389 10047
rect 29788 10016 30389 10044
rect 29788 10004 29794 10016
rect 30377 10013 30389 10016
rect 30423 10013 30435 10047
rect 30377 10007 30435 10013
rect 30470 10047 30528 10053
rect 30470 10013 30482 10047
rect 30516 10013 30528 10047
rect 30576 10044 30604 10152
rect 30842 10047 30900 10053
rect 30842 10044 30854 10047
rect 30576 10016 30854 10044
rect 30470 10007 30528 10013
rect 30842 10013 30854 10016
rect 30888 10013 30900 10047
rect 30842 10007 30900 10013
rect 25792 9948 29684 9976
rect 29917 9979 29975 9985
rect 25225 9939 25283 9945
rect 29917 9945 29929 9979
rect 29963 9976 29975 9979
rect 29963 9948 30512 9976
rect 29963 9945 29975 9948
rect 29917 9939 29975 9945
rect 30484 9920 30512 9948
rect 30650 9936 30656 9988
rect 30708 9936 30714 9988
rect 30742 9936 30748 9988
rect 30800 9936 30806 9988
rect 24397 9911 24455 9917
rect 24397 9877 24409 9911
rect 24443 9877 24455 9911
rect 24397 9871 24455 9877
rect 24670 9868 24676 9920
rect 24728 9908 24734 9920
rect 24857 9911 24915 9917
rect 24857 9908 24869 9911
rect 24728 9880 24869 9908
rect 24728 9868 24734 9880
rect 24857 9877 24869 9880
rect 24903 9877 24915 9911
rect 24857 9871 24915 9877
rect 29273 9911 29331 9917
rect 29273 9877 29285 9911
rect 29319 9908 29331 9911
rect 29454 9908 29460 9920
rect 29319 9880 29460 9908
rect 29319 9877 29331 9880
rect 29273 9871 29331 9877
rect 29454 9868 29460 9880
rect 29512 9868 29518 9920
rect 30006 9868 30012 9920
rect 30064 9868 30070 9920
rect 30466 9868 30472 9920
rect 30524 9868 30530 9920
rect 31018 9868 31024 9920
rect 31076 9868 31082 9920
rect 1104 9818 31832 9840
rect 1104 9766 4922 9818
rect 4974 9766 4986 9818
rect 5038 9766 5050 9818
rect 5102 9766 5114 9818
rect 5166 9766 5178 9818
rect 5230 9766 5242 9818
rect 5294 9766 10922 9818
rect 10974 9766 10986 9818
rect 11038 9766 11050 9818
rect 11102 9766 11114 9818
rect 11166 9766 11178 9818
rect 11230 9766 11242 9818
rect 11294 9766 16922 9818
rect 16974 9766 16986 9818
rect 17038 9766 17050 9818
rect 17102 9766 17114 9818
rect 17166 9766 17178 9818
rect 17230 9766 17242 9818
rect 17294 9766 22922 9818
rect 22974 9766 22986 9818
rect 23038 9766 23050 9818
rect 23102 9766 23114 9818
rect 23166 9766 23178 9818
rect 23230 9766 23242 9818
rect 23294 9766 28922 9818
rect 28974 9766 28986 9818
rect 29038 9766 29050 9818
rect 29102 9766 29114 9818
rect 29166 9766 29178 9818
rect 29230 9766 29242 9818
rect 29294 9766 31832 9818
rect 1104 9744 31832 9766
rect 7190 9664 7196 9716
rect 7248 9704 7254 9716
rect 7248 9676 8340 9704
rect 7248 9664 7254 9676
rect 8312 9636 8340 9676
rect 8386 9664 8392 9716
rect 8444 9664 8450 9716
rect 11238 9704 11244 9716
rect 8496 9676 11244 9704
rect 8496 9636 8524 9676
rect 11238 9664 11244 9676
rect 11296 9664 11302 9716
rect 11333 9707 11391 9713
rect 11333 9673 11345 9707
rect 11379 9673 11391 9707
rect 11333 9667 11391 9673
rect 8312 9608 8524 9636
rect 11348 9636 11376 9667
rect 12894 9664 12900 9716
rect 12952 9664 12958 9716
rect 18785 9707 18843 9713
rect 18785 9673 18797 9707
rect 18831 9673 18843 9707
rect 18785 9667 18843 9673
rect 11762 9639 11820 9645
rect 11762 9636 11774 9639
rect 11348 9608 11774 9636
rect 11762 9605 11774 9608
rect 11808 9605 11820 9639
rect 11762 9599 11820 9605
rect 2498 9528 2504 9580
rect 2556 9528 2562 9580
rect 2774 9577 2780 9580
rect 2768 9531 2780 9577
rect 2774 9528 2780 9531
rect 2832 9528 2838 9580
rect 7282 9577 7288 9580
rect 7276 9531 7288 9577
rect 7282 9528 7288 9531
rect 7340 9528 7346 9580
rect 11146 9528 11152 9580
rect 11204 9528 11210 9580
rect 11517 9571 11575 9577
rect 11517 9537 11529 9571
rect 11563 9568 11575 9571
rect 11606 9568 11612 9580
rect 11563 9540 11612 9568
rect 11563 9537 11575 9540
rect 11517 9531 11575 9537
rect 11606 9528 11612 9540
rect 11664 9528 11670 9580
rect 12912 9568 12940 9664
rect 14176 9639 14234 9645
rect 14176 9605 14188 9639
rect 14222 9636 14234 9639
rect 14642 9636 14648 9648
rect 14222 9608 14648 9636
rect 14222 9605 14234 9608
rect 14176 9599 14234 9605
rect 14642 9596 14648 9608
rect 14700 9596 14706 9648
rect 15746 9596 15752 9648
rect 15804 9636 15810 9648
rect 16117 9639 16175 9645
rect 16117 9636 16129 9639
rect 15804 9608 16129 9636
rect 15804 9596 15810 9608
rect 16117 9605 16129 9608
rect 16163 9605 16175 9639
rect 18800 9636 18828 9667
rect 20254 9664 20260 9716
rect 20312 9664 20318 9716
rect 20346 9664 20352 9716
rect 20404 9664 20410 9716
rect 21266 9664 21272 9716
rect 21324 9704 21330 9716
rect 23658 9704 23664 9716
rect 21324 9676 23664 9704
rect 21324 9664 21330 9676
rect 23658 9664 23664 9676
rect 23716 9664 23722 9716
rect 30006 9704 30012 9716
rect 28276 9676 30012 9704
rect 25130 9645 25136 9648
rect 19122 9639 19180 9645
rect 19122 9636 19134 9639
rect 18800 9608 19134 9636
rect 16117 9599 16175 9605
rect 19122 9605 19134 9608
rect 19168 9605 19180 9639
rect 20809 9639 20867 9645
rect 20809 9636 20821 9639
rect 19122 9599 19180 9605
rect 19444 9608 20821 9636
rect 19444 9580 19472 9608
rect 20809 9605 20821 9608
rect 20855 9605 20867 9639
rect 25102 9639 25136 9645
rect 20809 9599 20867 9605
rect 23400 9608 24900 9636
rect 13541 9571 13599 9577
rect 13541 9568 13553 9571
rect 12912 9540 13553 9568
rect 13541 9537 13553 9540
rect 13587 9537 13599 9571
rect 13541 9531 13599 9537
rect 13814 9528 13820 9580
rect 13872 9568 13878 9580
rect 13909 9571 13967 9577
rect 13909 9568 13921 9571
rect 13872 9540 13921 9568
rect 13872 9528 13878 9540
rect 13909 9537 13921 9540
rect 13955 9537 13967 9571
rect 13909 9531 13967 9537
rect 16301 9571 16359 9577
rect 16301 9537 16313 9571
rect 16347 9537 16359 9571
rect 16301 9531 16359 9537
rect 18601 9571 18659 9577
rect 18601 9537 18613 9571
rect 18647 9537 18659 9571
rect 18601 9531 18659 9537
rect 18877 9571 18935 9577
rect 18877 9537 18889 9571
rect 18923 9568 18935 9571
rect 18966 9568 18972 9580
rect 18923 9540 18972 9568
rect 18923 9537 18935 9540
rect 18877 9531 18935 9537
rect 6914 9460 6920 9512
rect 6972 9500 6978 9512
rect 7009 9503 7067 9509
rect 7009 9500 7021 9503
rect 6972 9472 7021 9500
rect 6972 9460 6978 9472
rect 7009 9469 7021 9472
rect 7055 9469 7067 9503
rect 15933 9503 15991 9509
rect 15933 9500 15945 9503
rect 7009 9463 7067 9469
rect 15304 9472 15945 9500
rect 3881 9435 3939 9441
rect 3881 9401 3893 9435
rect 3927 9432 3939 9435
rect 4706 9432 4712 9444
rect 3927 9404 4712 9432
rect 3927 9401 3939 9404
rect 3881 9395 3939 9401
rect 4706 9392 4712 9404
rect 4764 9392 4770 9444
rect 15304 9441 15332 9472
rect 15933 9469 15945 9472
rect 15979 9500 15991 9503
rect 16316 9500 16344 9531
rect 15979 9472 16344 9500
rect 15979 9469 15991 9472
rect 15933 9463 15991 9469
rect 15289 9435 15347 9441
rect 15289 9401 15301 9435
rect 15335 9401 15347 9435
rect 15289 9395 15347 9401
rect 12986 9324 12992 9376
rect 13044 9324 13050 9376
rect 15378 9324 15384 9376
rect 15436 9324 15442 9376
rect 15746 9324 15752 9376
rect 15804 9364 15810 9376
rect 16485 9367 16543 9373
rect 16485 9364 16497 9367
rect 15804 9336 16497 9364
rect 15804 9324 15810 9336
rect 16485 9333 16497 9336
rect 16531 9333 16543 9367
rect 18616 9364 18644 9531
rect 18966 9528 18972 9540
rect 19024 9528 19030 9580
rect 19426 9528 19432 9580
rect 19484 9528 19490 9580
rect 20714 9528 20720 9580
rect 20772 9528 20778 9580
rect 23106 9528 23112 9580
rect 23164 9528 23170 9580
rect 23400 9577 23428 9608
rect 24872 9577 24900 9608
rect 25102 9605 25114 9639
rect 25102 9599 25136 9605
rect 25130 9596 25136 9599
rect 25188 9596 25194 9648
rect 28074 9596 28080 9648
rect 28132 9636 28138 9648
rect 28276 9645 28304 9676
rect 30006 9664 30012 9676
rect 30064 9664 30070 9716
rect 30190 9664 30196 9716
rect 30248 9664 30254 9716
rect 30466 9664 30472 9716
rect 30524 9664 30530 9716
rect 28261 9639 28319 9645
rect 28261 9636 28273 9639
rect 28132 9608 28273 9636
rect 28132 9596 28138 9608
rect 28261 9605 28273 9608
rect 28307 9605 28319 9639
rect 28261 9599 28319 9605
rect 28353 9639 28411 9645
rect 28353 9605 28365 9639
rect 28399 9636 28411 9639
rect 28810 9636 28816 9648
rect 28399 9608 28816 9636
rect 28399 9605 28411 9608
rect 28353 9599 28411 9605
rect 28810 9596 28816 9608
rect 28868 9596 28874 9648
rect 29086 9645 29092 9648
rect 29080 9599 29092 9645
rect 29086 9596 29092 9599
rect 29144 9596 29150 9648
rect 29638 9596 29644 9648
rect 29696 9596 29702 9648
rect 23385 9571 23443 9577
rect 23385 9537 23397 9571
rect 23431 9537 23443 9571
rect 23641 9571 23699 9577
rect 23641 9568 23653 9571
rect 23385 9531 23443 9537
rect 23492 9540 23653 9568
rect 20993 9503 21051 9509
rect 20993 9469 21005 9503
rect 21039 9500 21051 9503
rect 23492 9500 23520 9540
rect 23641 9537 23653 9540
rect 23687 9537 23699 9571
rect 23641 9531 23699 9537
rect 24857 9571 24915 9577
rect 24857 9537 24869 9571
rect 24903 9568 24915 9571
rect 24946 9568 24952 9580
rect 24903 9540 24952 9568
rect 24903 9537 24915 9540
rect 24857 9531 24915 9537
rect 24946 9528 24952 9540
rect 25004 9528 25010 9580
rect 25682 9528 25688 9580
rect 25740 9568 25746 9580
rect 29656 9568 29684 9596
rect 25740 9540 29684 9568
rect 25740 9528 25746 9540
rect 28184 9509 28212 9540
rect 30742 9528 30748 9580
rect 30800 9568 30806 9580
rect 31021 9571 31079 9577
rect 31021 9568 31033 9571
rect 30800 9540 31033 9568
rect 30800 9528 30806 9540
rect 31021 9537 31033 9540
rect 31067 9537 31079 9571
rect 31021 9531 31079 9537
rect 21039 9472 22094 9500
rect 21039 9469 21051 9472
rect 20993 9463 21051 9469
rect 19242 9364 19248 9376
rect 18616 9336 19248 9364
rect 16485 9327 16543 9333
rect 19242 9324 19248 9336
rect 19300 9324 19306 9376
rect 22066 9364 22094 9472
rect 23308 9472 23520 9500
rect 28169 9503 28227 9509
rect 23308 9441 23336 9472
rect 28169 9469 28181 9503
rect 28215 9469 28227 9503
rect 28169 9463 28227 9469
rect 28810 9460 28816 9512
rect 28868 9509 28874 9512
rect 28868 9500 28878 9509
rect 28868 9472 28913 9500
rect 28868 9463 28878 9472
rect 28868 9460 28874 9463
rect 23293 9435 23351 9441
rect 23293 9401 23305 9435
rect 23339 9401 23351 9435
rect 23293 9395 23351 9401
rect 24486 9364 24492 9376
rect 22066 9336 24492 9364
rect 24486 9324 24492 9336
rect 24544 9324 24550 9376
rect 24762 9324 24768 9376
rect 24820 9324 24826 9376
rect 26050 9324 26056 9376
rect 26108 9364 26114 9376
rect 26237 9367 26295 9373
rect 26237 9364 26249 9367
rect 26108 9336 26249 9364
rect 26108 9324 26114 9336
rect 26237 9333 26249 9336
rect 26283 9333 26295 9367
rect 26237 9327 26295 9333
rect 28718 9324 28724 9376
rect 28776 9324 28782 9376
rect 1104 9274 31832 9296
rect 1104 9222 4182 9274
rect 4234 9222 4246 9274
rect 4298 9222 4310 9274
rect 4362 9222 4374 9274
rect 4426 9222 4438 9274
rect 4490 9222 4502 9274
rect 4554 9222 10182 9274
rect 10234 9222 10246 9274
rect 10298 9222 10310 9274
rect 10362 9222 10374 9274
rect 10426 9222 10438 9274
rect 10490 9222 10502 9274
rect 10554 9222 16182 9274
rect 16234 9222 16246 9274
rect 16298 9222 16310 9274
rect 16362 9222 16374 9274
rect 16426 9222 16438 9274
rect 16490 9222 16502 9274
rect 16554 9222 22182 9274
rect 22234 9222 22246 9274
rect 22298 9222 22310 9274
rect 22362 9222 22374 9274
rect 22426 9222 22438 9274
rect 22490 9222 22502 9274
rect 22554 9222 28182 9274
rect 28234 9222 28246 9274
rect 28298 9222 28310 9274
rect 28362 9222 28374 9274
rect 28426 9222 28438 9274
rect 28490 9222 28502 9274
rect 28554 9222 31832 9274
rect 1104 9200 31832 9222
rect 2774 9120 2780 9172
rect 2832 9160 2838 9172
rect 2869 9163 2927 9169
rect 2869 9160 2881 9163
rect 2832 9132 2881 9160
rect 2832 9120 2838 9132
rect 2869 9129 2881 9132
rect 2915 9129 2927 9163
rect 2869 9123 2927 9129
rect 7282 9120 7288 9172
rect 7340 9160 7346 9172
rect 7469 9163 7527 9169
rect 7469 9160 7481 9163
rect 7340 9132 7481 9160
rect 7340 9120 7346 9132
rect 7469 9129 7481 9132
rect 7515 9129 7527 9163
rect 7469 9123 7527 9129
rect 11146 9120 11152 9172
rect 11204 9160 11210 9172
rect 11885 9163 11943 9169
rect 11885 9160 11897 9163
rect 11204 9132 11897 9160
rect 11204 9120 11210 9132
rect 11885 9129 11897 9132
rect 11931 9129 11943 9163
rect 11885 9123 11943 9129
rect 14826 9120 14832 9172
rect 14884 9160 14890 9172
rect 15105 9163 15163 9169
rect 15105 9160 15117 9163
rect 14884 9132 15117 9160
rect 14884 9120 14890 9132
rect 15105 9129 15117 9132
rect 15151 9129 15163 9163
rect 15105 9123 15163 9129
rect 15378 9120 15384 9172
rect 15436 9120 15442 9172
rect 18506 9120 18512 9172
rect 18564 9120 18570 9172
rect 19061 9163 19119 9169
rect 19061 9129 19073 9163
rect 19107 9160 19119 9163
rect 19702 9160 19708 9172
rect 19107 9132 19708 9160
rect 19107 9129 19119 9132
rect 19061 9123 19119 9129
rect 19702 9120 19708 9132
rect 19760 9120 19766 9172
rect 20714 9120 20720 9172
rect 20772 9160 20778 9172
rect 20809 9163 20867 9169
rect 20809 9160 20821 9163
rect 20772 9132 20821 9160
rect 20772 9120 20778 9132
rect 20809 9129 20821 9132
rect 20855 9129 20867 9163
rect 20809 9123 20867 9129
rect 22830 9120 22836 9172
rect 22888 9120 22894 9172
rect 23106 9120 23112 9172
rect 23164 9160 23170 9172
rect 24397 9163 24455 9169
rect 24397 9160 24409 9163
rect 23164 9132 24409 9160
rect 23164 9120 23170 9132
rect 24397 9129 24409 9132
rect 24443 9129 24455 9163
rect 26050 9160 26056 9172
rect 24397 9123 24455 9129
rect 24688 9132 26056 9160
rect 8754 9052 8760 9104
rect 8812 9052 8818 9104
rect 11241 9095 11299 9101
rect 11241 9061 11253 9095
rect 11287 9092 11299 9095
rect 11330 9092 11336 9104
rect 11287 9064 11336 9092
rect 11287 9061 11299 9064
rect 11241 9055 11299 9061
rect 11330 9052 11336 9064
rect 11388 9052 11394 9104
rect 8772 9024 8800 9052
rect 11149 9027 11207 9033
rect 11149 9024 11161 9027
rect 8772 8996 11161 9024
rect 11149 8993 11161 8996
rect 11195 8993 11207 9027
rect 11149 8987 11207 8993
rect 12158 8984 12164 9036
rect 12216 9024 12222 9036
rect 12529 9027 12587 9033
rect 12529 9024 12541 9027
rect 12216 8996 12541 9024
rect 12216 8984 12222 8996
rect 12529 8993 12541 8996
rect 12575 9024 12587 9027
rect 14553 9027 14611 9033
rect 14553 9024 14565 9027
rect 12575 8996 14565 9024
rect 12575 8993 12587 8996
rect 12529 8987 12587 8993
rect 14553 8993 14565 8996
rect 14599 9024 14611 9027
rect 15010 9024 15016 9036
rect 14599 8996 15016 9024
rect 14599 8993 14611 8996
rect 14553 8987 14611 8993
rect 15010 8984 15016 8996
rect 15068 8984 15074 9036
rect 3053 8959 3111 8965
rect 3053 8925 3065 8959
rect 3099 8956 3111 8959
rect 3786 8956 3792 8968
rect 3099 8928 3792 8956
rect 3099 8925 3111 8928
rect 3053 8919 3111 8925
rect 3786 8916 3792 8928
rect 3844 8916 3850 8968
rect 7653 8959 7711 8965
rect 7653 8925 7665 8959
rect 7699 8956 7711 8959
rect 7926 8956 7932 8968
rect 7699 8928 7932 8956
rect 7699 8925 7711 8928
rect 7653 8919 7711 8925
rect 7926 8916 7932 8928
rect 7984 8916 7990 8968
rect 9766 8916 9772 8968
rect 9824 8956 9830 8968
rect 10137 8959 10195 8965
rect 10137 8956 10149 8959
rect 9824 8928 10149 8956
rect 9824 8916 9830 8928
rect 10137 8925 10149 8928
rect 10183 8925 10195 8959
rect 10137 8919 10195 8925
rect 11057 8959 11115 8965
rect 11057 8925 11069 8959
rect 11103 8925 11115 8959
rect 11057 8919 11115 8925
rect 11333 8959 11391 8965
rect 11333 8925 11345 8959
rect 11379 8956 11391 8959
rect 11514 8956 11520 8968
rect 11379 8928 11520 8956
rect 11379 8925 11391 8928
rect 11333 8919 11391 8925
rect 10686 8848 10692 8900
rect 10744 8888 10750 8900
rect 10873 8891 10931 8897
rect 10873 8888 10885 8891
rect 10744 8860 10885 8888
rect 10744 8848 10750 8860
rect 10873 8857 10885 8860
rect 10919 8857 10931 8891
rect 11072 8888 11100 8919
rect 11514 8916 11520 8928
rect 11572 8916 11578 8968
rect 12253 8959 12311 8965
rect 12253 8925 12265 8959
rect 12299 8956 12311 8959
rect 12986 8956 12992 8968
rect 12299 8928 12992 8956
rect 12299 8925 12311 8928
rect 12253 8919 12311 8925
rect 12986 8916 12992 8928
rect 13044 8916 13050 8968
rect 14737 8959 14795 8965
rect 14737 8925 14749 8959
rect 14783 8956 14795 8959
rect 15396 8956 15424 9120
rect 18524 9092 18552 9120
rect 19334 9092 19340 9104
rect 18524 9064 19340 9092
rect 17589 9027 17647 9033
rect 17589 8993 17601 9027
rect 17635 9024 17647 9027
rect 18524 9024 18552 9064
rect 19334 9052 19340 9064
rect 19392 9052 19398 9104
rect 23017 9095 23075 9101
rect 23017 9092 23029 9095
rect 20364 9064 23029 9092
rect 17635 8996 18552 9024
rect 17635 8993 17647 8996
rect 17589 8987 17647 8993
rect 18325 8959 18383 8965
rect 14783 8928 15424 8956
rect 17236 8928 17908 8956
rect 14783 8925 14795 8928
rect 14737 8919 14795 8925
rect 17236 8888 17264 8928
rect 11072 8860 17264 8888
rect 17313 8891 17371 8897
rect 10873 8851 10931 8857
rect 17313 8857 17325 8891
rect 17359 8888 17371 8891
rect 17773 8891 17831 8897
rect 17773 8888 17785 8891
rect 17359 8860 17785 8888
rect 17359 8857 17371 8860
rect 17313 8851 17371 8857
rect 17773 8857 17785 8860
rect 17819 8857 17831 8891
rect 17773 8851 17831 8857
rect 8570 8780 8576 8832
rect 8628 8820 8634 8832
rect 10318 8820 10324 8832
rect 8628 8792 10324 8820
rect 8628 8780 8634 8792
rect 10318 8780 10324 8792
rect 10376 8780 10382 8832
rect 10778 8780 10784 8832
rect 10836 8780 10842 8832
rect 12345 8823 12403 8829
rect 12345 8789 12357 8823
rect 12391 8820 12403 8823
rect 12434 8820 12440 8832
rect 12391 8792 12440 8820
rect 12391 8789 12403 8792
rect 12345 8783 12403 8789
rect 12434 8780 12440 8792
rect 12492 8780 12498 8832
rect 13814 8780 13820 8832
rect 13872 8820 13878 8832
rect 14366 8820 14372 8832
rect 13872 8792 14372 8820
rect 13872 8780 13878 8792
rect 14366 8780 14372 8792
rect 14424 8780 14430 8832
rect 14645 8823 14703 8829
rect 14645 8789 14657 8823
rect 14691 8820 14703 8823
rect 15102 8820 15108 8832
rect 14691 8792 15108 8820
rect 14691 8789 14703 8792
rect 14645 8783 14703 8789
rect 15102 8780 15108 8792
rect 15160 8780 15166 8832
rect 16482 8780 16488 8832
rect 16540 8820 16546 8832
rect 16945 8823 17003 8829
rect 16945 8820 16957 8823
rect 16540 8792 16957 8820
rect 16540 8780 16546 8792
rect 16945 8789 16957 8792
rect 16991 8789 17003 8823
rect 16945 8783 17003 8789
rect 17405 8823 17463 8829
rect 17405 8789 17417 8823
rect 17451 8820 17463 8823
rect 17678 8820 17684 8832
rect 17451 8792 17684 8820
rect 17451 8789 17463 8792
rect 17405 8783 17463 8789
rect 17678 8780 17684 8792
rect 17736 8780 17742 8832
rect 17880 8820 17908 8928
rect 18325 8925 18337 8959
rect 18371 8925 18383 8959
rect 18325 8919 18383 8925
rect 18046 8848 18052 8900
rect 18104 8888 18110 8900
rect 18340 8888 18368 8919
rect 18506 8916 18512 8968
rect 18564 8916 18570 8968
rect 18785 8959 18843 8965
rect 18785 8956 18797 8959
rect 18616 8928 18797 8956
rect 18616 8888 18644 8928
rect 18785 8925 18797 8928
rect 18831 8925 18843 8959
rect 18785 8919 18843 8925
rect 18877 8959 18935 8965
rect 18877 8925 18889 8959
rect 18923 8925 18935 8959
rect 18877 8919 18935 8925
rect 18104 8860 18644 8888
rect 18104 8848 18110 8860
rect 18690 8848 18696 8900
rect 18748 8848 18754 8900
rect 18892 8888 18920 8919
rect 18966 8916 18972 8968
rect 19024 8956 19030 8968
rect 19337 8959 19395 8965
rect 19337 8956 19349 8959
rect 19024 8928 19349 8956
rect 19024 8916 19030 8928
rect 19337 8925 19349 8928
rect 19383 8956 19395 8959
rect 19886 8956 19892 8968
rect 19383 8928 19892 8956
rect 19383 8925 19395 8928
rect 19337 8919 19395 8925
rect 19886 8916 19892 8928
rect 19944 8916 19950 8968
rect 20162 8916 20168 8968
rect 20220 8916 20226 8968
rect 19426 8888 19432 8900
rect 18892 8860 19432 8888
rect 19426 8848 19432 8860
rect 19484 8848 19490 8900
rect 19604 8891 19662 8897
rect 19604 8857 19616 8891
rect 19650 8888 19662 8891
rect 20180 8888 20208 8916
rect 19650 8860 20208 8888
rect 19650 8857 19662 8860
rect 19604 8851 19662 8857
rect 20364 8820 20392 9064
rect 23017 9061 23029 9064
rect 23063 9061 23075 9095
rect 24688 9092 24716 9132
rect 26050 9120 26056 9132
rect 26108 9120 26114 9172
rect 26418 9120 26424 9172
rect 26476 9120 26482 9172
rect 28718 9120 28724 9172
rect 28776 9120 28782 9172
rect 29086 9120 29092 9172
rect 29144 9160 29150 9172
rect 29181 9163 29239 9169
rect 29181 9160 29193 9163
rect 29144 9132 29193 9160
rect 29144 9120 29150 9132
rect 29181 9129 29193 9132
rect 29227 9129 29239 9163
rect 29181 9123 29239 9129
rect 30742 9120 30748 9172
rect 30800 9160 30806 9172
rect 30929 9163 30987 9169
rect 30929 9160 30941 9163
rect 30800 9132 30941 9160
rect 30800 9120 30806 9132
rect 30929 9129 30941 9132
rect 30975 9129 30987 9163
rect 30929 9123 30987 9129
rect 23017 9055 23075 9061
rect 23860 9064 24716 9092
rect 21174 8984 21180 9036
rect 21232 9024 21238 9036
rect 21361 9027 21419 9033
rect 21361 9024 21373 9027
rect 21232 8996 21373 9024
rect 21232 8984 21238 8996
rect 21361 8993 21373 8996
rect 21407 8993 21419 9027
rect 21361 8987 21419 8993
rect 21818 8984 21824 9036
rect 21876 9024 21882 9036
rect 22646 9024 22652 9036
rect 21876 8996 22652 9024
rect 21876 8984 21882 8996
rect 22646 8984 22652 8996
rect 22704 8984 22710 9036
rect 17880 8792 20392 8820
rect 20717 8823 20775 8829
rect 20717 8789 20729 8823
rect 20763 8820 20775 8823
rect 21192 8820 21220 8984
rect 22738 8916 22744 8968
rect 22796 8916 22802 8968
rect 23750 8965 23756 8968
rect 22833 8959 22891 8965
rect 22833 8925 22845 8959
rect 22879 8956 22891 8959
rect 23748 8956 23756 8965
rect 22879 8928 23612 8956
rect 23711 8928 23756 8956
rect 22879 8925 22891 8928
rect 22833 8919 22891 8925
rect 22557 8891 22615 8897
rect 22557 8857 22569 8891
rect 22603 8888 22615 8891
rect 22646 8888 22652 8900
rect 22603 8860 22652 8888
rect 22603 8857 22615 8860
rect 22557 8851 22615 8857
rect 22646 8848 22652 8860
rect 22704 8848 22710 8900
rect 20763 8792 21220 8820
rect 20763 8789 20775 8792
rect 20717 8783 20775 8789
rect 22094 8780 22100 8832
rect 22152 8820 22158 8832
rect 22830 8820 22836 8832
rect 22152 8792 22836 8820
rect 22152 8780 22158 8792
rect 22830 8780 22836 8792
rect 22888 8780 22894 8832
rect 23584 8829 23612 8928
rect 23748 8919 23756 8928
rect 23750 8916 23756 8919
rect 23808 8916 23814 8968
rect 23860 8965 23888 9064
rect 24762 9052 24768 9104
rect 24820 9092 24826 9104
rect 24820 9064 25820 9092
rect 24820 9052 24826 9064
rect 24780 9024 24808 9052
rect 24136 8996 24808 9024
rect 25041 9027 25099 9033
rect 24136 8965 24164 8996
rect 25041 8993 25053 9027
rect 25087 9024 25099 9027
rect 25682 9024 25688 9036
rect 25087 8996 25688 9024
rect 25087 8993 25099 8996
rect 25041 8987 25099 8993
rect 23845 8959 23903 8965
rect 23845 8925 23857 8959
rect 23891 8925 23903 8959
rect 23845 8919 23903 8925
rect 24120 8959 24178 8965
rect 24120 8925 24132 8959
rect 24166 8925 24178 8959
rect 24120 8919 24178 8925
rect 24213 8959 24271 8965
rect 24213 8925 24225 8959
rect 24259 8956 24271 8959
rect 24394 8956 24400 8968
rect 24259 8928 24400 8956
rect 24259 8925 24271 8928
rect 24213 8919 24271 8925
rect 24394 8916 24400 8928
rect 24452 8916 24458 8968
rect 24578 8916 24584 8968
rect 24636 8956 24642 8968
rect 25056 8956 25084 8987
rect 25682 8984 25688 8996
rect 25740 8984 25746 9036
rect 25792 9033 25820 9064
rect 25777 9027 25835 9033
rect 25777 8993 25789 9027
rect 25823 8993 25835 9027
rect 25777 8987 25835 8993
rect 24636 8928 25084 8956
rect 24636 8916 24642 8928
rect 26602 8916 26608 8968
rect 26660 8916 26666 8968
rect 26697 8959 26755 8965
rect 26697 8925 26709 8959
rect 26743 8925 26755 8959
rect 28736 8956 28764 9120
rect 28810 8984 28816 9036
rect 28868 9024 28874 9036
rect 29549 9027 29607 9033
rect 29549 9024 29561 9027
rect 28868 8996 29561 9024
rect 28868 8984 28874 8996
rect 29549 8993 29561 8996
rect 29595 8993 29607 9027
rect 29549 8987 29607 8993
rect 28997 8959 29055 8965
rect 28997 8956 29009 8959
rect 28736 8928 29009 8956
rect 26697 8919 26755 8925
rect 28997 8925 29009 8928
rect 29043 8925 29055 8959
rect 28997 8919 29055 8925
rect 23937 8891 23995 8897
rect 23937 8857 23949 8891
rect 23983 8857 23995 8891
rect 23937 8851 23995 8857
rect 24765 8891 24823 8897
rect 24765 8857 24777 8891
rect 24811 8888 24823 8891
rect 25225 8891 25283 8897
rect 25225 8888 25237 8891
rect 24811 8860 25237 8888
rect 24811 8857 24823 8860
rect 24765 8851 24823 8857
rect 25225 8857 25237 8860
rect 25271 8857 25283 8891
rect 25225 8851 25283 8857
rect 23569 8823 23627 8829
rect 23569 8789 23581 8823
rect 23615 8789 23627 8823
rect 23569 8783 23627 8789
rect 23658 8780 23664 8832
rect 23716 8820 23722 8832
rect 23952 8820 23980 8851
rect 26418 8848 26424 8900
rect 26476 8848 26482 8900
rect 26712 8888 26740 8919
rect 29454 8916 29460 8968
rect 29512 8956 29518 8968
rect 29805 8959 29863 8965
rect 29805 8956 29817 8959
rect 29512 8928 29817 8956
rect 29512 8916 29518 8928
rect 29805 8925 29817 8928
rect 29851 8925 29863 8959
rect 29805 8919 29863 8925
rect 31018 8916 31024 8968
rect 31076 8916 31082 8968
rect 31036 8888 31064 8916
rect 26712 8860 31064 8888
rect 23716 8792 23980 8820
rect 23716 8780 23722 8792
rect 24854 8780 24860 8832
rect 24912 8780 24918 8832
rect 26878 8780 26884 8832
rect 26936 8780 26942 8832
rect 1104 8730 31832 8752
rect 1104 8678 4922 8730
rect 4974 8678 4986 8730
rect 5038 8678 5050 8730
rect 5102 8678 5114 8730
rect 5166 8678 5178 8730
rect 5230 8678 5242 8730
rect 5294 8678 10922 8730
rect 10974 8678 10986 8730
rect 11038 8678 11050 8730
rect 11102 8678 11114 8730
rect 11166 8678 11178 8730
rect 11230 8678 11242 8730
rect 11294 8678 16922 8730
rect 16974 8678 16986 8730
rect 17038 8678 17050 8730
rect 17102 8678 17114 8730
rect 17166 8678 17178 8730
rect 17230 8678 17242 8730
rect 17294 8678 22922 8730
rect 22974 8678 22986 8730
rect 23038 8678 23050 8730
rect 23102 8678 23114 8730
rect 23166 8678 23178 8730
rect 23230 8678 23242 8730
rect 23294 8678 28922 8730
rect 28974 8678 28986 8730
rect 29038 8678 29050 8730
rect 29102 8678 29114 8730
rect 29166 8678 29178 8730
rect 29230 8678 29242 8730
rect 29294 8678 31832 8730
rect 1104 8656 31832 8678
rect 9858 8576 9864 8628
rect 9916 8576 9922 8628
rect 10505 8619 10563 8625
rect 10505 8585 10517 8619
rect 10551 8616 10563 8619
rect 10778 8616 10784 8628
rect 10551 8588 10784 8616
rect 10551 8585 10563 8588
rect 10505 8579 10563 8585
rect 10778 8576 10784 8588
rect 10836 8576 10842 8628
rect 13814 8616 13820 8628
rect 12406 8588 13820 8616
rect 9585 8551 9643 8557
rect 7392 8520 9352 8548
rect 5994 8440 6000 8492
rect 6052 8440 6058 8492
rect 6638 8372 6644 8424
rect 6696 8412 6702 8424
rect 7392 8421 7420 8520
rect 8113 8483 8171 8489
rect 8113 8449 8125 8483
rect 8159 8449 8171 8483
rect 8113 8443 8171 8449
rect 8297 8483 8355 8489
rect 8297 8449 8309 8483
rect 8343 8449 8355 8483
rect 8297 8443 8355 8449
rect 7377 8415 7435 8421
rect 7377 8412 7389 8415
rect 6696 8384 7389 8412
rect 6696 8372 6702 8384
rect 7377 8381 7389 8384
rect 7423 8381 7435 8415
rect 7377 8375 7435 8381
rect 5810 8304 5816 8356
rect 5868 8304 5874 8356
rect 8128 8344 8156 8443
rect 8312 8412 8340 8443
rect 8386 8440 8392 8492
rect 8444 8440 8450 8492
rect 8481 8483 8539 8489
rect 8481 8449 8493 8483
rect 8527 8480 8539 8483
rect 8938 8480 8944 8492
rect 8527 8452 8944 8480
rect 8527 8449 8539 8452
rect 8481 8443 8539 8449
rect 8938 8440 8944 8452
rect 8996 8440 9002 8492
rect 9214 8440 9220 8492
rect 9272 8440 9278 8492
rect 9324 8489 9352 8520
rect 9585 8517 9597 8551
rect 9631 8548 9643 8551
rect 9950 8548 9956 8560
rect 9631 8520 9956 8548
rect 9631 8517 9643 8520
rect 9585 8511 9643 8517
rect 9950 8508 9956 8520
rect 10008 8508 10014 8560
rect 12406 8548 12434 8588
rect 13814 8576 13820 8588
rect 13872 8576 13878 8628
rect 13998 8576 14004 8628
rect 14056 8616 14062 8628
rect 14056 8588 14228 8616
rect 14056 8576 14062 8588
rect 14200 8557 14228 8588
rect 15746 8576 15752 8628
rect 15804 8576 15810 8628
rect 16482 8576 16488 8628
rect 16540 8576 16546 8628
rect 18046 8576 18052 8628
rect 18104 8576 18110 8628
rect 18141 8619 18199 8625
rect 18141 8585 18153 8619
rect 18187 8585 18199 8619
rect 19150 8616 19156 8628
rect 18141 8579 18199 8585
rect 18432 8588 19156 8616
rect 10520 8520 12434 8548
rect 14185 8551 14243 8557
rect 9310 8483 9368 8489
rect 9310 8449 9322 8483
rect 9356 8449 9368 8483
rect 9310 8443 9368 8449
rect 9493 8483 9551 8489
rect 9493 8449 9505 8483
rect 9539 8449 9551 8483
rect 9493 8443 9551 8449
rect 9508 8412 9536 8443
rect 9674 8440 9680 8492
rect 9732 8489 9738 8492
rect 9732 8483 9781 8489
rect 9732 8449 9735 8483
rect 9769 8480 9781 8483
rect 10520 8480 10548 8520
rect 14185 8517 14197 8551
rect 14231 8517 14243 8551
rect 14185 8511 14243 8517
rect 14277 8551 14335 8557
rect 14277 8517 14289 8551
rect 14323 8548 14335 8551
rect 15470 8548 15476 8560
rect 14323 8520 15476 8548
rect 14323 8517 14335 8520
rect 14277 8511 14335 8517
rect 12434 8480 12440 8492
rect 9769 8452 10548 8480
rect 10612 8452 12440 8480
rect 9769 8449 9781 8452
rect 9732 8443 9781 8449
rect 9732 8440 9738 8443
rect 8312 8384 8524 8412
rect 8496 8356 8524 8384
rect 9508 8384 10272 8412
rect 8294 8344 8300 8356
rect 8128 8316 8300 8344
rect 8294 8304 8300 8316
rect 8352 8304 8358 8356
rect 8478 8304 8484 8356
rect 8536 8304 8542 8356
rect 9306 8304 9312 8356
rect 9364 8344 9370 8356
rect 9508 8344 9536 8384
rect 9364 8316 9536 8344
rect 9364 8304 9370 8316
rect 10042 8304 10048 8356
rect 10100 8344 10106 8356
rect 10137 8347 10195 8353
rect 10137 8344 10149 8347
rect 10100 8316 10149 8344
rect 10100 8304 10106 8316
rect 10137 8313 10149 8316
rect 10183 8313 10195 8347
rect 10244 8344 10272 8384
rect 10318 8372 10324 8424
rect 10376 8412 10382 8424
rect 10612 8421 10640 8452
rect 12434 8440 12440 8452
rect 12492 8440 12498 8492
rect 13722 8440 13728 8492
rect 13780 8480 13786 8492
rect 14090 8489 14096 8492
rect 13909 8483 13967 8489
rect 13909 8480 13921 8483
rect 13780 8452 13921 8480
rect 13780 8440 13786 8452
rect 13909 8449 13921 8452
rect 13955 8449 13967 8483
rect 13909 8443 13967 8449
rect 14057 8483 14096 8489
rect 14057 8449 14069 8483
rect 14057 8443 14096 8449
rect 14090 8440 14096 8443
rect 14148 8440 14154 8492
rect 10597 8415 10655 8421
rect 10597 8412 10609 8415
rect 10376 8384 10609 8412
rect 10376 8372 10382 8384
rect 10597 8381 10609 8384
rect 10643 8381 10655 8415
rect 10597 8375 10655 8381
rect 10778 8372 10784 8424
rect 10836 8372 10842 8424
rect 14200 8344 14228 8511
rect 15470 8508 15476 8520
rect 15528 8508 15534 8560
rect 14366 8440 14372 8492
rect 14424 8489 14430 8492
rect 14424 8480 14432 8489
rect 14424 8452 14469 8480
rect 14424 8443 14432 8452
rect 14424 8440 14430 8443
rect 14550 8440 14556 8492
rect 14608 8480 14614 8492
rect 14645 8483 14703 8489
rect 14645 8480 14657 8483
rect 14608 8452 14657 8480
rect 14608 8440 14614 8452
rect 14645 8449 14657 8452
rect 14691 8449 14703 8483
rect 14645 8443 14703 8449
rect 14826 8440 14832 8492
rect 14884 8440 14890 8492
rect 14918 8440 14924 8492
rect 14976 8440 14982 8492
rect 15105 8483 15163 8489
rect 15105 8449 15117 8483
rect 15151 8480 15163 8483
rect 15764 8480 15792 8576
rect 16500 8548 16528 8576
rect 18156 8548 18184 8579
rect 16040 8520 16528 8548
rect 16592 8520 18184 8548
rect 16040 8489 16068 8520
rect 15151 8452 15792 8480
rect 16025 8483 16083 8489
rect 15151 8449 15163 8452
rect 15105 8443 15163 8449
rect 16025 8449 16037 8483
rect 16071 8449 16083 8483
rect 16025 8443 16083 8449
rect 16301 8483 16359 8489
rect 16301 8449 16313 8483
rect 16347 8480 16359 8483
rect 16592 8480 16620 8520
rect 16347 8452 16620 8480
rect 16347 8449 16359 8452
rect 16301 8443 16359 8449
rect 16666 8440 16672 8492
rect 16724 8440 16730 8492
rect 16925 8483 16983 8489
rect 16925 8480 16937 8483
rect 16776 8452 16937 8480
rect 15013 8415 15071 8421
rect 15013 8412 15025 8415
rect 14568 8384 15025 8412
rect 14568 8353 14596 8384
rect 15013 8381 15025 8384
rect 15059 8381 15071 8415
rect 16776 8412 16804 8452
rect 16925 8449 16937 8452
rect 16971 8449 16983 8483
rect 16925 8443 16983 8449
rect 18432 8412 18460 8588
rect 19150 8576 19156 8588
rect 19208 8576 19214 8628
rect 19426 8576 19432 8628
rect 19484 8616 19490 8628
rect 20438 8616 20444 8628
rect 19484 8588 20444 8616
rect 19484 8576 19490 8588
rect 20438 8576 20444 8588
rect 20496 8616 20502 8628
rect 22465 8619 22523 8625
rect 20496 8588 22324 8616
rect 20496 8576 20502 8588
rect 18690 8508 18696 8560
rect 18748 8548 18754 8560
rect 19978 8548 19984 8560
rect 18748 8520 19984 8548
rect 18748 8508 18754 8520
rect 19978 8508 19984 8520
rect 20036 8548 20042 8560
rect 22094 8548 22100 8560
rect 20036 8520 22100 8548
rect 20036 8508 20042 8520
rect 22094 8508 22100 8520
rect 22152 8508 22158 8560
rect 18509 8483 18567 8489
rect 18509 8449 18521 8483
rect 18555 8480 18567 8483
rect 18969 8483 19027 8489
rect 18969 8480 18981 8483
rect 18555 8452 18981 8480
rect 18555 8449 18567 8452
rect 18509 8443 18567 8449
rect 18969 8449 18981 8452
rect 19015 8449 19027 8483
rect 18969 8443 19027 8449
rect 21913 8483 21971 8489
rect 21913 8449 21925 8483
rect 21959 8480 21971 8483
rect 21959 8452 22094 8480
rect 21959 8449 21971 8452
rect 21913 8443 21971 8449
rect 18601 8415 18659 8421
rect 18601 8412 18613 8415
rect 15013 8375 15071 8381
rect 16224 8384 16804 8412
rect 17696 8384 18613 8412
rect 16224 8353 16252 8384
rect 10244 8316 14228 8344
rect 14553 8347 14611 8353
rect 10137 8307 10195 8313
rect 14553 8313 14565 8347
rect 14599 8313 14611 8347
rect 14553 8307 14611 8313
rect 16209 8347 16267 8353
rect 16209 8313 16221 8347
rect 16255 8313 16267 8347
rect 16209 8307 16267 8313
rect 16485 8347 16543 8353
rect 16485 8313 16497 8347
rect 16531 8344 16543 8347
rect 16531 8316 16712 8344
rect 16531 8313 16543 8316
rect 16485 8307 16543 8313
rect 6546 8236 6552 8288
rect 6604 8276 6610 8288
rect 6825 8279 6883 8285
rect 6825 8276 6837 8279
rect 6604 8248 6837 8276
rect 6604 8236 6610 8248
rect 6825 8245 6837 8248
rect 6871 8245 6883 8279
rect 6825 8239 6883 8245
rect 8662 8236 8668 8288
rect 8720 8236 8726 8288
rect 9858 8236 9864 8288
rect 9916 8276 9922 8288
rect 10778 8276 10784 8288
rect 9916 8248 10784 8276
rect 9916 8236 9922 8248
rect 10778 8236 10784 8248
rect 10836 8236 10842 8288
rect 16684 8276 16712 8316
rect 16850 8276 16856 8288
rect 16684 8248 16856 8276
rect 16850 8236 16856 8248
rect 16908 8236 16914 8288
rect 17310 8236 17316 8288
rect 17368 8276 17374 8288
rect 17696 8276 17724 8384
rect 18601 8381 18613 8384
rect 18647 8381 18659 8415
rect 18601 8375 18659 8381
rect 18785 8415 18843 8421
rect 18785 8381 18797 8415
rect 18831 8412 18843 8415
rect 19426 8412 19432 8424
rect 18831 8384 19432 8412
rect 18831 8381 18843 8384
rect 18785 8375 18843 8381
rect 19426 8372 19432 8384
rect 19484 8372 19490 8424
rect 19521 8415 19579 8421
rect 19521 8381 19533 8415
rect 19567 8381 19579 8415
rect 22066 8412 22094 8452
rect 22186 8440 22192 8492
rect 22244 8440 22250 8492
rect 22296 8489 22324 8588
rect 22465 8585 22477 8619
rect 22511 8616 22523 8619
rect 22738 8616 22744 8628
rect 22511 8588 22744 8616
rect 22511 8585 22523 8588
rect 22465 8579 22523 8585
rect 22738 8576 22744 8588
rect 22796 8576 22802 8628
rect 26237 8619 26295 8625
rect 26237 8585 26249 8619
rect 26283 8616 26295 8619
rect 26602 8616 26608 8628
rect 26283 8588 26608 8616
rect 26283 8585 26295 8588
rect 26237 8579 26295 8585
rect 26602 8576 26608 8588
rect 26660 8576 26666 8628
rect 27338 8616 27344 8628
rect 26804 8588 27344 8616
rect 22830 8508 22836 8560
rect 22888 8548 22894 8560
rect 22888 8520 26648 8548
rect 22888 8508 22894 8520
rect 26620 8489 26648 8520
rect 26804 8489 26832 8588
rect 27338 8576 27344 8588
rect 27396 8576 27402 8628
rect 27080 8520 28488 8548
rect 22281 8483 22339 8489
rect 22281 8449 22293 8483
rect 22327 8480 22339 8483
rect 26421 8483 26479 8489
rect 26421 8480 26433 8483
rect 22327 8452 26433 8480
rect 22327 8449 22339 8452
rect 22281 8443 22339 8449
rect 26421 8449 26433 8452
rect 26467 8449 26479 8483
rect 26421 8443 26479 8449
rect 26513 8483 26571 8489
rect 26513 8449 26525 8483
rect 26559 8449 26571 8483
rect 26513 8443 26571 8449
rect 26605 8483 26663 8489
rect 26605 8449 26617 8483
rect 26651 8449 26663 8483
rect 26605 8443 26663 8449
rect 26789 8483 26847 8489
rect 26789 8449 26801 8483
rect 26835 8449 26847 8483
rect 26789 8443 26847 8449
rect 23382 8412 23388 8424
rect 22066 8384 23388 8412
rect 19521 8375 19579 8381
rect 18506 8304 18512 8356
rect 18564 8344 18570 8356
rect 19536 8344 19564 8375
rect 23382 8372 23388 8384
rect 23440 8372 23446 8424
rect 26528 8412 26556 8443
rect 27080 8424 27108 8520
rect 28460 8489 28488 8520
rect 27433 8483 27491 8489
rect 27433 8449 27445 8483
rect 27479 8480 27491 8483
rect 27893 8483 27951 8489
rect 27893 8480 27905 8483
rect 27479 8452 27905 8480
rect 27479 8449 27491 8452
rect 27433 8443 27491 8449
rect 27893 8449 27905 8452
rect 27939 8449 27951 8483
rect 27893 8443 27951 8449
rect 28445 8483 28503 8489
rect 28445 8449 28457 8483
rect 28491 8449 28503 8483
rect 28445 8443 28503 8449
rect 28629 8483 28687 8489
rect 28629 8449 28641 8483
rect 28675 8480 28687 8483
rect 29362 8480 29368 8492
rect 28675 8452 29368 8480
rect 28675 8449 28687 8452
rect 28629 8443 28687 8449
rect 27062 8412 27068 8424
rect 26528 8384 27068 8412
rect 27062 8372 27068 8384
rect 27120 8372 27126 8424
rect 27157 8415 27215 8421
rect 27157 8381 27169 8415
rect 27203 8381 27215 8415
rect 27157 8375 27215 8381
rect 27341 8415 27399 8421
rect 27341 8381 27353 8415
rect 27387 8412 27399 8415
rect 28644 8412 28672 8443
rect 29362 8440 29368 8452
rect 29420 8440 29426 8492
rect 27387 8384 28672 8412
rect 27387 8381 27399 8384
rect 27341 8375 27399 8381
rect 18564 8316 19564 8344
rect 18564 8304 18570 8316
rect 22738 8304 22744 8356
rect 22796 8344 22802 8356
rect 27172 8344 27200 8375
rect 22796 8316 27200 8344
rect 22796 8304 22802 8316
rect 17368 8248 17724 8276
rect 17368 8236 17374 8248
rect 24670 8236 24676 8288
rect 24728 8276 24734 8288
rect 27356 8276 27384 8375
rect 28074 8344 28080 8356
rect 27448 8316 28080 8344
rect 27448 8288 27476 8316
rect 28074 8304 28080 8316
rect 28132 8344 28138 8356
rect 28813 8347 28871 8353
rect 28813 8344 28825 8347
rect 28132 8316 28825 8344
rect 28132 8304 28138 8316
rect 28813 8313 28825 8316
rect 28859 8313 28871 8347
rect 28813 8307 28871 8313
rect 24728 8248 27384 8276
rect 24728 8236 24734 8248
rect 27430 8236 27436 8288
rect 27488 8236 27494 8288
rect 27798 8236 27804 8288
rect 27856 8236 27862 8288
rect 1104 8186 31832 8208
rect 1104 8134 4182 8186
rect 4234 8134 4246 8186
rect 4298 8134 4310 8186
rect 4362 8134 4374 8186
rect 4426 8134 4438 8186
rect 4490 8134 4502 8186
rect 4554 8134 10182 8186
rect 10234 8134 10246 8186
rect 10298 8134 10310 8186
rect 10362 8134 10374 8186
rect 10426 8134 10438 8186
rect 10490 8134 10502 8186
rect 10554 8134 16182 8186
rect 16234 8134 16246 8186
rect 16298 8134 16310 8186
rect 16362 8134 16374 8186
rect 16426 8134 16438 8186
rect 16490 8134 16502 8186
rect 16554 8134 22182 8186
rect 22234 8134 22246 8186
rect 22298 8134 22310 8186
rect 22362 8134 22374 8186
rect 22426 8134 22438 8186
rect 22490 8134 22502 8186
rect 22554 8134 28182 8186
rect 28234 8134 28246 8186
rect 28298 8134 28310 8186
rect 28362 8134 28374 8186
rect 28426 8134 28438 8186
rect 28490 8134 28502 8186
rect 28554 8134 31832 8186
rect 1104 8112 31832 8134
rect 9766 8072 9772 8084
rect 9416 8044 9772 8072
rect 6641 8007 6699 8013
rect 6641 7973 6653 8007
rect 6687 8004 6699 8007
rect 6687 7976 8156 8004
rect 6687 7973 6699 7976
rect 6641 7967 6699 7973
rect 2498 7896 2504 7948
rect 2556 7936 2562 7948
rect 8128 7945 8156 7976
rect 5261 7939 5319 7945
rect 5261 7936 5273 7939
rect 2556 7908 5273 7936
rect 2556 7896 2562 7908
rect 5261 7905 5273 7908
rect 5307 7905 5319 7939
rect 5261 7899 5319 7905
rect 7377 7939 7435 7945
rect 7377 7905 7389 7939
rect 7423 7905 7435 7939
rect 7377 7899 7435 7905
rect 8113 7939 8171 7945
rect 8113 7905 8125 7939
rect 8159 7936 8171 7939
rect 8159 7908 9168 7936
rect 8159 7905 8171 7908
rect 8113 7899 8171 7905
rect 5276 7868 5304 7899
rect 5350 7868 5356 7880
rect 5276 7840 5356 7868
rect 5350 7828 5356 7840
rect 5408 7828 5414 7880
rect 7282 7828 7288 7880
rect 7340 7868 7346 7880
rect 7392 7868 7420 7899
rect 7340 7840 7420 7868
rect 7340 7828 7346 7840
rect 8662 7828 8668 7880
rect 8720 7868 8726 7880
rect 9140 7877 9168 7908
rect 9033 7871 9091 7877
rect 9033 7868 9045 7871
rect 8720 7840 9045 7868
rect 8720 7828 8726 7840
rect 9033 7837 9045 7840
rect 9079 7837 9091 7871
rect 9033 7831 9091 7837
rect 9126 7871 9184 7877
rect 9126 7837 9138 7871
rect 9172 7837 9184 7871
rect 9126 7831 9184 7837
rect 9306 7828 9312 7880
rect 9364 7828 9370 7880
rect 9416 7877 9444 8044
rect 9766 8032 9772 8044
rect 9824 8032 9830 8084
rect 17957 8075 18015 8081
rect 17957 8041 17969 8075
rect 18003 8072 18015 8075
rect 18506 8072 18512 8084
rect 18003 8044 18512 8072
rect 18003 8041 18015 8044
rect 17957 8035 18015 8041
rect 18506 8032 18512 8044
rect 18564 8032 18570 8084
rect 19334 8032 19340 8084
rect 19392 8072 19398 8084
rect 20622 8072 20628 8084
rect 19392 8044 20628 8072
rect 19392 8032 19398 8044
rect 20622 8032 20628 8044
rect 20680 8072 20686 8084
rect 22738 8072 22744 8084
rect 20680 8044 22744 8072
rect 20680 8032 20686 8044
rect 22738 8032 22744 8044
rect 22796 8032 22802 8084
rect 27062 8032 27068 8084
rect 27120 8072 27126 8084
rect 27525 8075 27583 8081
rect 27525 8072 27537 8075
rect 27120 8044 27537 8072
rect 27120 8032 27126 8044
rect 27525 8041 27537 8044
rect 27571 8041 27583 8075
rect 27525 8035 27583 8041
rect 31110 8032 31116 8084
rect 31168 8032 31174 8084
rect 13354 8004 13360 8016
rect 12544 7976 13360 8004
rect 12544 7948 12572 7976
rect 13354 7964 13360 7976
rect 13412 8004 13418 8016
rect 13412 7976 14688 8004
rect 13412 7964 13418 7976
rect 11149 7939 11207 7945
rect 11149 7905 11161 7939
rect 11195 7936 11207 7939
rect 11606 7936 11612 7948
rect 11195 7908 11612 7936
rect 11195 7905 11207 7908
rect 11149 7899 11207 7905
rect 11606 7896 11612 7908
rect 11664 7896 11670 7948
rect 12526 7896 12532 7948
rect 12584 7896 12590 7948
rect 13464 7908 13676 7936
rect 9401 7871 9459 7877
rect 9401 7837 9413 7871
rect 9447 7837 9459 7871
rect 9401 7831 9459 7837
rect 9539 7871 9597 7877
rect 9539 7837 9551 7871
rect 9585 7868 9597 7871
rect 9674 7868 9680 7880
rect 9585 7840 9680 7868
rect 9585 7837 9597 7840
rect 9539 7831 9597 7837
rect 9674 7828 9680 7840
rect 9732 7828 9738 7880
rect 11330 7828 11336 7880
rect 11388 7828 11394 7880
rect 5528 7803 5586 7809
rect 5528 7769 5540 7803
rect 5574 7800 5586 7803
rect 5626 7800 5632 7812
rect 5574 7772 5632 7800
rect 5574 7769 5586 7772
rect 5528 7763 5586 7769
rect 5626 7760 5632 7772
rect 5684 7760 5690 7812
rect 7101 7803 7159 7809
rect 7101 7769 7113 7803
rect 7147 7800 7159 7803
rect 7561 7803 7619 7809
rect 7561 7800 7573 7803
rect 7147 7772 7573 7800
rect 7147 7769 7159 7772
rect 7101 7763 7159 7769
rect 7561 7769 7573 7772
rect 7607 7769 7619 7803
rect 7561 7763 7619 7769
rect 9766 7760 9772 7812
rect 9824 7800 9830 7812
rect 10502 7800 10508 7812
rect 9824 7772 10508 7800
rect 9824 7760 9830 7772
rect 10502 7760 10508 7772
rect 10560 7760 10566 7812
rect 10686 7760 10692 7812
rect 10744 7800 10750 7812
rect 10882 7803 10940 7809
rect 10882 7800 10894 7803
rect 10744 7772 10894 7800
rect 10744 7760 10750 7772
rect 10882 7769 10894 7772
rect 10928 7769 10940 7803
rect 10882 7763 10940 7769
rect 6730 7692 6736 7744
rect 6788 7692 6794 7744
rect 7193 7735 7251 7741
rect 7193 7701 7205 7735
rect 7239 7732 7251 7735
rect 7466 7732 7472 7744
rect 7239 7704 7472 7732
rect 7239 7701 7251 7704
rect 7193 7695 7251 7701
rect 7466 7692 7472 7704
rect 7524 7692 7530 7744
rect 9677 7735 9735 7741
rect 9677 7701 9689 7735
rect 9723 7732 9735 7735
rect 11348 7732 11376 7828
rect 11422 7760 11428 7812
rect 11480 7800 11486 7812
rect 12250 7800 12256 7812
rect 11480 7772 12256 7800
rect 11480 7760 11486 7772
rect 12250 7760 12256 7772
rect 12308 7800 12314 7812
rect 13464 7800 13492 7908
rect 13541 7871 13599 7877
rect 13541 7837 13553 7871
rect 13587 7837 13599 7871
rect 13541 7831 13599 7837
rect 12308 7772 13492 7800
rect 12308 7760 12314 7772
rect 9723 7704 11376 7732
rect 13357 7735 13415 7741
rect 9723 7701 9735 7704
rect 9677 7695 9735 7701
rect 13357 7701 13369 7735
rect 13403 7732 13415 7735
rect 13446 7732 13452 7744
rect 13403 7704 13452 7732
rect 13403 7701 13415 7704
rect 13357 7695 13415 7701
rect 13446 7692 13452 7704
rect 13504 7692 13510 7744
rect 13556 7732 13584 7831
rect 13648 7800 13676 7908
rect 14090 7896 14096 7948
rect 14148 7936 14154 7948
rect 14660 7945 14688 7976
rect 19426 7964 19432 8016
rect 19484 8004 19490 8016
rect 19794 8004 19800 8016
rect 19484 7976 19800 8004
rect 19484 7964 19490 7976
rect 19794 7964 19800 7976
rect 19852 8004 19858 8016
rect 19852 7976 22600 8004
rect 19852 7964 19858 7976
rect 14645 7939 14703 7945
rect 14148 7908 14596 7936
rect 14148 7896 14154 7908
rect 14568 7868 14596 7908
rect 14645 7905 14657 7939
rect 14691 7905 14703 7939
rect 14645 7899 14703 7905
rect 20622 7896 20628 7948
rect 20680 7896 20686 7948
rect 21545 7939 21603 7945
rect 21545 7905 21557 7939
rect 21591 7936 21603 7939
rect 22094 7936 22100 7948
rect 21591 7908 22100 7936
rect 21591 7905 21603 7908
rect 21545 7899 21603 7905
rect 22094 7896 22100 7908
rect 22152 7896 22158 7948
rect 22572 7945 22600 7976
rect 22557 7939 22615 7945
rect 22557 7905 22569 7939
rect 22603 7936 22615 7939
rect 22830 7936 22836 7948
rect 22603 7908 22836 7936
rect 22603 7905 22615 7908
rect 22557 7899 22615 7905
rect 22830 7896 22836 7908
rect 22888 7896 22894 7948
rect 23382 7896 23388 7948
rect 23440 7896 23446 7948
rect 24854 7896 24860 7948
rect 24912 7896 24918 7948
rect 15473 7871 15531 7877
rect 15473 7868 15485 7871
rect 14568 7840 15485 7868
rect 15473 7837 15485 7840
rect 15519 7837 15531 7871
rect 15473 7831 15531 7837
rect 16577 7871 16635 7877
rect 16577 7837 16589 7871
rect 16623 7868 16635 7871
rect 16666 7868 16672 7880
rect 16623 7840 16672 7868
rect 16623 7837 16635 7840
rect 16577 7831 16635 7837
rect 16666 7828 16672 7840
rect 16724 7828 16730 7880
rect 16850 7877 16856 7880
rect 16844 7868 16856 7877
rect 16811 7840 16856 7868
rect 16844 7831 16856 7840
rect 16850 7828 16856 7831
rect 16908 7828 16914 7880
rect 21818 7828 21824 7880
rect 21876 7868 21882 7880
rect 22373 7871 22431 7877
rect 22373 7868 22385 7871
rect 21876 7840 22385 7868
rect 21876 7828 21882 7840
rect 22373 7837 22385 7840
rect 22419 7868 22431 7871
rect 24872 7868 24900 7896
rect 22419 7840 24900 7868
rect 22419 7837 22431 7840
rect 22373 7831 22431 7837
rect 25774 7828 25780 7880
rect 25832 7828 25838 7880
rect 26053 7871 26111 7877
rect 26053 7868 26065 7871
rect 25884 7840 26065 7868
rect 14461 7803 14519 7809
rect 13648 7772 14412 7800
rect 14093 7735 14151 7741
rect 14093 7732 14105 7735
rect 13556 7704 14105 7732
rect 14093 7701 14105 7704
rect 14139 7701 14151 7735
rect 14384 7732 14412 7772
rect 14461 7769 14473 7803
rect 14507 7800 14519 7803
rect 14921 7803 14979 7809
rect 14921 7800 14933 7803
rect 14507 7772 14933 7800
rect 14507 7769 14519 7772
rect 14461 7763 14519 7769
rect 14921 7769 14933 7772
rect 14967 7769 14979 7803
rect 14921 7763 14979 7769
rect 20441 7803 20499 7809
rect 20441 7769 20453 7803
rect 20487 7800 20499 7803
rect 20901 7803 20959 7809
rect 20901 7800 20913 7803
rect 20487 7772 20913 7800
rect 20487 7769 20499 7772
rect 20441 7763 20499 7769
rect 20901 7769 20913 7772
rect 20947 7769 20959 7803
rect 20901 7763 20959 7769
rect 22281 7803 22339 7809
rect 22281 7769 22293 7803
rect 22327 7800 22339 7803
rect 22833 7803 22891 7809
rect 22833 7800 22845 7803
rect 22327 7772 22845 7800
rect 22327 7769 22339 7772
rect 22281 7763 22339 7769
rect 22833 7769 22845 7772
rect 22879 7769 22891 7803
rect 22833 7763 22891 7769
rect 23658 7760 23664 7812
rect 23716 7800 23722 7812
rect 24946 7800 24952 7812
rect 23716 7772 24952 7800
rect 23716 7760 23722 7772
rect 24946 7760 24952 7772
rect 25004 7800 25010 7812
rect 25884 7800 25912 7840
rect 26053 7837 26065 7840
rect 26099 7868 26111 7871
rect 28810 7868 28816 7880
rect 26099 7840 28816 7868
rect 26099 7837 26111 7840
rect 26053 7831 26111 7837
rect 28810 7828 28816 7840
rect 28868 7868 28874 7880
rect 28905 7871 28963 7877
rect 28905 7868 28917 7871
rect 28868 7840 28917 7868
rect 28868 7828 28874 7840
rect 28905 7837 28917 7840
rect 28951 7837 28963 7871
rect 28905 7831 28963 7837
rect 26298 7803 26356 7809
rect 26298 7800 26310 7803
rect 25004 7772 25912 7800
rect 25976 7772 26310 7800
rect 25004 7760 25010 7772
rect 14553 7735 14611 7741
rect 14553 7732 14565 7735
rect 14384 7704 14565 7732
rect 14093 7695 14151 7701
rect 14553 7701 14565 7704
rect 14599 7732 14611 7735
rect 16574 7732 16580 7744
rect 14599 7704 16580 7732
rect 14599 7701 14611 7704
rect 14553 7695 14611 7701
rect 16574 7692 16580 7704
rect 16632 7692 16638 7744
rect 19610 7692 19616 7744
rect 19668 7732 19674 7744
rect 20073 7735 20131 7741
rect 20073 7732 20085 7735
rect 19668 7704 20085 7732
rect 19668 7692 19674 7704
rect 20073 7701 20085 7704
rect 20119 7701 20131 7735
rect 20073 7695 20131 7701
rect 20533 7735 20591 7741
rect 20533 7701 20545 7735
rect 20579 7732 20591 7735
rect 20622 7732 20628 7744
rect 20579 7704 20628 7732
rect 20579 7701 20591 7704
rect 20533 7695 20591 7701
rect 20622 7692 20628 7704
rect 20680 7692 20686 7744
rect 21634 7692 21640 7744
rect 21692 7732 21698 7744
rect 25976 7741 26004 7772
rect 26298 7769 26310 7772
rect 26344 7769 26356 7803
rect 26298 7763 26356 7769
rect 28626 7760 28632 7812
rect 28684 7809 28690 7812
rect 28684 7763 28696 7809
rect 31389 7803 31447 7809
rect 31389 7769 31401 7803
rect 31435 7800 31447 7803
rect 31846 7800 31852 7812
rect 31435 7772 31852 7800
rect 31435 7769 31447 7772
rect 31389 7763 31447 7769
rect 28684 7760 28690 7763
rect 31846 7760 31852 7772
rect 31904 7760 31910 7812
rect 21913 7735 21971 7741
rect 21913 7732 21925 7735
rect 21692 7704 21925 7732
rect 21692 7692 21698 7704
rect 21913 7701 21925 7704
rect 21959 7701 21971 7735
rect 21913 7695 21971 7701
rect 25961 7735 26019 7741
rect 25961 7701 25973 7735
rect 26007 7701 26019 7735
rect 25961 7695 26019 7701
rect 27338 7692 27344 7744
rect 27396 7732 27402 7744
rect 27433 7735 27491 7741
rect 27433 7732 27445 7735
rect 27396 7704 27445 7732
rect 27396 7692 27402 7704
rect 27433 7701 27445 7704
rect 27479 7701 27491 7735
rect 27433 7695 27491 7701
rect 1104 7642 31832 7664
rect 1104 7590 4922 7642
rect 4974 7590 4986 7642
rect 5038 7590 5050 7642
rect 5102 7590 5114 7642
rect 5166 7590 5178 7642
rect 5230 7590 5242 7642
rect 5294 7590 10922 7642
rect 10974 7590 10986 7642
rect 11038 7590 11050 7642
rect 11102 7590 11114 7642
rect 11166 7590 11178 7642
rect 11230 7590 11242 7642
rect 11294 7590 16922 7642
rect 16974 7590 16986 7642
rect 17038 7590 17050 7642
rect 17102 7590 17114 7642
rect 17166 7590 17178 7642
rect 17230 7590 17242 7642
rect 17294 7590 22922 7642
rect 22974 7590 22986 7642
rect 23038 7590 23050 7642
rect 23102 7590 23114 7642
rect 23166 7590 23178 7642
rect 23230 7590 23242 7642
rect 23294 7590 28922 7642
rect 28974 7590 28986 7642
rect 29038 7590 29050 7642
rect 29102 7590 29114 7642
rect 29166 7590 29178 7642
rect 29230 7590 29242 7642
rect 29294 7590 31832 7642
rect 1104 7568 31832 7590
rect 5626 7488 5632 7540
rect 5684 7488 5690 7540
rect 5994 7488 6000 7540
rect 6052 7528 6058 7540
rect 6365 7531 6423 7537
rect 6365 7528 6377 7531
rect 6052 7500 6377 7528
rect 6052 7488 6058 7500
rect 6365 7497 6377 7500
rect 6411 7497 6423 7531
rect 6365 7491 6423 7497
rect 6546 7488 6552 7540
rect 6604 7528 6610 7540
rect 6733 7531 6791 7537
rect 6733 7528 6745 7531
rect 6604 7500 6745 7528
rect 6604 7488 6610 7500
rect 6733 7497 6745 7500
rect 6779 7497 6791 7531
rect 6733 7491 6791 7497
rect 6825 7531 6883 7537
rect 6825 7497 6837 7531
rect 6871 7528 6883 7531
rect 7653 7531 7711 7537
rect 7653 7528 7665 7531
rect 6871 7500 7665 7528
rect 6871 7497 6883 7500
rect 6825 7491 6883 7497
rect 7653 7497 7665 7500
rect 7699 7528 7711 7531
rect 7699 7500 9168 7528
rect 7699 7497 7711 7500
rect 7653 7491 7711 7497
rect 5902 7420 5908 7472
rect 5960 7460 5966 7472
rect 6840 7460 6868 7491
rect 5960 7432 6868 7460
rect 5960 7420 5966 7432
rect 6914 7420 6920 7472
rect 6972 7460 6978 7472
rect 8846 7460 8852 7472
rect 6972 7432 8852 7460
rect 6972 7420 6978 7432
rect 8846 7420 8852 7432
rect 8904 7420 8910 7472
rect 9140 7460 9168 7500
rect 9950 7488 9956 7540
rect 10008 7528 10014 7540
rect 10413 7531 10471 7537
rect 10413 7528 10425 7531
rect 10008 7500 10425 7528
rect 10008 7488 10014 7500
rect 10413 7497 10425 7500
rect 10459 7497 10471 7531
rect 10413 7491 10471 7497
rect 9674 7460 9680 7472
rect 9140 7432 9680 7460
rect 9674 7420 9680 7432
rect 9732 7420 9738 7472
rect 10428 7460 10456 7491
rect 10502 7488 10508 7540
rect 10560 7528 10566 7540
rect 10560 7500 13308 7528
rect 10560 7488 10566 7500
rect 13280 7460 13308 7500
rect 14090 7488 14096 7540
rect 14148 7528 14154 7540
rect 14553 7531 14611 7537
rect 14553 7528 14565 7531
rect 14148 7500 14565 7528
rect 14148 7488 14154 7500
rect 14553 7497 14565 7500
rect 14599 7497 14611 7531
rect 14553 7491 14611 7497
rect 19610 7488 19616 7540
rect 19668 7488 19674 7540
rect 21637 7531 21695 7537
rect 19904 7500 21588 7528
rect 10428 7432 11100 7460
rect 13280 7432 14780 7460
rect 5813 7395 5871 7401
rect 5813 7361 5825 7395
rect 5859 7392 5871 7395
rect 6730 7392 6736 7404
rect 5859 7364 6736 7392
rect 5859 7361 5871 7364
rect 5813 7355 5871 7361
rect 6730 7352 6736 7364
rect 6788 7352 6794 7404
rect 7561 7395 7619 7401
rect 7561 7361 7573 7395
rect 7607 7392 7619 7395
rect 8021 7395 8079 7401
rect 8021 7392 8033 7395
rect 7607 7364 8033 7392
rect 7607 7361 7619 7364
rect 7561 7355 7619 7361
rect 8021 7361 8033 7364
rect 8067 7361 8079 7395
rect 8021 7355 8079 7361
rect 8754 7352 8760 7404
rect 8812 7352 8818 7404
rect 8864 7392 8892 7420
rect 11072 7401 11100 7432
rect 9022 7395 9080 7401
rect 9022 7392 9034 7395
rect 8864 7364 9034 7392
rect 9022 7361 9034 7364
rect 9068 7361 9080 7395
rect 9289 7395 9347 7401
rect 9289 7392 9301 7395
rect 9022 7355 9080 7361
rect 9140 7364 9301 7392
rect 7009 7327 7067 7333
rect 7009 7293 7021 7327
rect 7055 7324 7067 7327
rect 7282 7324 7288 7336
rect 7055 7296 7288 7324
rect 7055 7293 7067 7296
rect 7009 7287 7067 7293
rect 7282 7284 7288 7296
rect 7340 7284 7346 7336
rect 7742 7284 7748 7336
rect 7800 7324 7806 7336
rect 7837 7327 7895 7333
rect 7837 7324 7849 7327
rect 7800 7296 7849 7324
rect 7800 7284 7806 7296
rect 7837 7293 7849 7296
rect 7883 7324 7895 7327
rect 8202 7324 8208 7336
rect 7883 7296 8208 7324
rect 7883 7293 7895 7296
rect 7837 7287 7895 7293
rect 8202 7284 8208 7296
rect 8260 7284 8266 7336
rect 8570 7284 8576 7336
rect 8628 7284 8634 7336
rect 9140 7324 9168 7364
rect 9289 7361 9301 7364
rect 9335 7361 9347 7395
rect 9289 7355 9347 7361
rect 11057 7395 11115 7401
rect 11057 7361 11069 7395
rect 11103 7361 11115 7395
rect 11057 7355 11115 7361
rect 11606 7352 11612 7404
rect 11664 7392 11670 7404
rect 13446 7401 13452 7404
rect 13429 7395 13452 7401
rect 11664 7364 13216 7392
rect 11664 7352 11670 7364
rect 12526 7324 12532 7336
rect 8956 7296 9168 7324
rect 10060 7296 12532 7324
rect 7190 7148 7196 7200
rect 7248 7148 7254 7200
rect 7300 7188 7328 7284
rect 8956 7265 8984 7296
rect 8941 7259 8999 7265
rect 8941 7225 8953 7259
rect 8987 7225 8999 7259
rect 8941 7219 8999 7225
rect 10060 7188 10088 7296
rect 12526 7284 12532 7296
rect 12584 7284 12590 7336
rect 13188 7333 13216 7364
rect 13429 7361 13441 7395
rect 13429 7355 13452 7361
rect 13446 7352 13452 7355
rect 13504 7352 13510 7404
rect 14752 7336 14780 7432
rect 15013 7395 15071 7401
rect 15013 7361 15025 7395
rect 15059 7392 15071 7395
rect 15473 7395 15531 7401
rect 15473 7392 15485 7395
rect 15059 7364 15485 7392
rect 15059 7361 15071 7364
rect 15013 7355 15071 7361
rect 15473 7361 15485 7364
rect 15519 7361 15531 7395
rect 15473 7355 15531 7361
rect 19521 7395 19579 7401
rect 19521 7361 19533 7395
rect 19567 7392 19579 7395
rect 19628 7392 19656 7488
rect 19904 7472 19932 7500
rect 19886 7460 19892 7472
rect 19812 7432 19892 7460
rect 19812 7401 19840 7432
rect 19886 7420 19892 7432
rect 19944 7420 19950 7472
rect 21560 7460 21588 7500
rect 21637 7497 21649 7531
rect 21683 7528 21695 7531
rect 23201 7531 23259 7537
rect 21683 7500 22094 7528
rect 21683 7497 21695 7500
rect 21637 7491 21695 7497
rect 22066 7469 22094 7500
rect 23201 7497 23213 7531
rect 23247 7528 23259 7531
rect 23382 7528 23388 7540
rect 23247 7500 23388 7528
rect 23247 7497 23259 7500
rect 23201 7491 23259 7497
rect 23382 7488 23388 7500
rect 23440 7488 23446 7540
rect 25774 7488 25780 7540
rect 25832 7528 25838 7540
rect 26973 7531 27031 7537
rect 26973 7528 26985 7531
rect 25832 7500 26985 7528
rect 25832 7488 25838 7500
rect 26973 7497 26985 7500
rect 27019 7497 27031 7531
rect 26973 7491 27031 7497
rect 27798 7488 27804 7540
rect 27856 7488 27862 7540
rect 28626 7488 28632 7540
rect 28684 7528 28690 7540
rect 28721 7531 28779 7537
rect 28721 7528 28733 7531
rect 28684 7500 28733 7528
rect 28684 7488 28690 7500
rect 28721 7497 28733 7500
rect 28767 7497 28779 7531
rect 28721 7491 28779 7497
rect 22066 7463 22124 7469
rect 21560 7432 21864 7460
rect 19567 7364 19656 7392
rect 19797 7395 19855 7401
rect 19567 7361 19579 7364
rect 19521 7355 19579 7361
rect 19797 7361 19809 7395
rect 19843 7361 19855 7395
rect 20053 7395 20111 7401
rect 20053 7392 20065 7395
rect 19797 7355 19855 7361
rect 19904 7364 20065 7392
rect 13173 7327 13231 7333
rect 13173 7293 13185 7327
rect 13219 7293 13231 7327
rect 13173 7287 13231 7293
rect 7300 7160 10088 7188
rect 10505 7191 10563 7197
rect 10505 7157 10517 7191
rect 10551 7188 10563 7191
rect 10870 7188 10876 7200
rect 10551 7160 10876 7188
rect 10551 7157 10563 7160
rect 10505 7151 10563 7157
rect 10870 7148 10876 7160
rect 10928 7148 10934 7200
rect 13188 7188 13216 7287
rect 14734 7284 14740 7336
rect 14792 7284 14798 7336
rect 15102 7284 15108 7336
rect 15160 7284 15166 7336
rect 15197 7327 15255 7333
rect 15197 7293 15209 7327
rect 15243 7293 15255 7327
rect 16025 7327 16083 7333
rect 16025 7324 16037 7327
rect 15197 7287 15255 7293
rect 15488 7296 16037 7324
rect 14752 7256 14780 7284
rect 15212 7256 15240 7287
rect 15488 7268 15516 7296
rect 16025 7293 16037 7296
rect 16071 7293 16083 7327
rect 19904 7324 19932 7364
rect 20053 7361 20065 7364
rect 20099 7361 20111 7395
rect 20053 7355 20111 7361
rect 21453 7395 21511 7401
rect 21453 7361 21465 7395
rect 21499 7392 21511 7395
rect 21634 7392 21640 7404
rect 21499 7364 21640 7392
rect 21499 7361 21511 7364
rect 21453 7355 21511 7361
rect 21634 7352 21640 7364
rect 21692 7352 21698 7404
rect 21836 7401 21864 7432
rect 22066 7429 22078 7463
rect 22112 7429 22124 7463
rect 27430 7460 27436 7472
rect 22066 7423 22124 7429
rect 25608 7432 27436 7460
rect 25608 7404 25636 7432
rect 27430 7420 27436 7432
rect 27488 7420 27494 7472
rect 21821 7395 21879 7401
rect 21821 7361 21833 7395
rect 21867 7361 21879 7395
rect 21821 7355 21879 7361
rect 25590 7352 25596 7404
rect 25648 7352 25654 7404
rect 27341 7395 27399 7401
rect 27341 7361 27353 7395
rect 27387 7392 27399 7395
rect 27816 7392 27844 7488
rect 28537 7395 28595 7401
rect 28537 7392 28549 7395
rect 27387 7364 27660 7392
rect 27816 7364 28549 7392
rect 27387 7361 27399 7364
rect 27341 7355 27399 7361
rect 16025 7287 16083 7293
rect 19720 7296 19932 7324
rect 14752 7228 15240 7256
rect 15470 7216 15476 7268
rect 15528 7216 15534 7268
rect 19720 7265 19748 7296
rect 22830 7284 22836 7336
rect 22888 7324 22894 7336
rect 27525 7327 27583 7333
rect 27525 7324 27537 7327
rect 22888 7296 27537 7324
rect 22888 7284 22894 7296
rect 27525 7293 27537 7296
rect 27571 7293 27583 7327
rect 27632 7324 27660 7364
rect 28537 7361 28549 7364
rect 28583 7361 28595 7395
rect 28537 7355 28595 7361
rect 27801 7327 27859 7333
rect 27801 7324 27813 7327
rect 27632 7296 27813 7324
rect 27525 7287 27583 7293
rect 27801 7293 27813 7296
rect 27847 7293 27859 7327
rect 27801 7287 27859 7293
rect 28353 7327 28411 7333
rect 28353 7293 28365 7327
rect 28399 7293 28411 7327
rect 28353 7287 28411 7293
rect 19705 7259 19763 7265
rect 19705 7225 19717 7259
rect 19751 7225 19763 7259
rect 19705 7219 19763 7225
rect 21192 7228 21772 7256
rect 13446 7188 13452 7200
rect 13188 7160 13452 7188
rect 13446 7148 13452 7160
rect 13504 7148 13510 7200
rect 14642 7148 14648 7200
rect 14700 7148 14706 7200
rect 21192 7197 21220 7228
rect 21177 7191 21235 7197
rect 21177 7157 21189 7191
rect 21223 7157 21235 7191
rect 21744 7188 21772 7228
rect 27338 7216 27344 7268
rect 27396 7256 27402 7268
rect 28368 7256 28396 7287
rect 27396 7228 28396 7256
rect 27396 7216 27402 7228
rect 22094 7188 22100 7200
rect 21744 7160 22100 7188
rect 21177 7151 21235 7157
rect 22094 7148 22100 7160
rect 22152 7148 22158 7200
rect 1104 7098 31832 7120
rect 1104 7046 4182 7098
rect 4234 7046 4246 7098
rect 4298 7046 4310 7098
rect 4362 7046 4374 7098
rect 4426 7046 4438 7098
rect 4490 7046 4502 7098
rect 4554 7046 10182 7098
rect 10234 7046 10246 7098
rect 10298 7046 10310 7098
rect 10362 7046 10374 7098
rect 10426 7046 10438 7098
rect 10490 7046 10502 7098
rect 10554 7046 16182 7098
rect 16234 7046 16246 7098
rect 16298 7046 16310 7098
rect 16362 7046 16374 7098
rect 16426 7046 16438 7098
rect 16490 7046 16502 7098
rect 16554 7046 22182 7098
rect 22234 7046 22246 7098
rect 22298 7046 22310 7098
rect 22362 7046 22374 7098
rect 22426 7046 22438 7098
rect 22490 7046 22502 7098
rect 22554 7046 28182 7098
rect 28234 7046 28246 7098
rect 28298 7046 28310 7098
rect 28362 7046 28374 7098
rect 28426 7046 28438 7098
rect 28490 7046 28502 7098
rect 28554 7046 31832 7098
rect 1104 7024 31832 7046
rect 8754 6944 8760 6996
rect 8812 6984 8818 6996
rect 9493 6987 9551 6993
rect 9493 6984 9505 6987
rect 8812 6956 9505 6984
rect 8812 6944 8818 6956
rect 9493 6953 9505 6956
rect 9539 6953 9551 6987
rect 9493 6947 9551 6953
rect 10686 6944 10692 6996
rect 10744 6944 10750 6996
rect 12066 6944 12072 6996
rect 12124 6944 12130 6996
rect 15378 6944 15384 6996
rect 15436 6944 15442 6996
rect 15470 6944 15476 6996
rect 15528 6944 15534 6996
rect 16574 6944 16580 6996
rect 16632 6984 16638 6996
rect 24670 6984 24676 6996
rect 16632 6956 24676 6984
rect 16632 6944 16638 6956
rect 24670 6944 24676 6956
rect 24728 6944 24734 6996
rect 8202 6876 8208 6928
rect 8260 6916 8266 6928
rect 12084 6916 12112 6944
rect 8260 6888 12112 6916
rect 8260 6876 8266 6888
rect 13722 6876 13728 6928
rect 13780 6876 13786 6928
rect 15396 6916 15424 6944
rect 15396 6888 17172 6916
rect 5350 6808 5356 6860
rect 5408 6848 5414 6860
rect 5445 6851 5503 6857
rect 5445 6848 5457 6851
rect 5408 6820 5457 6848
rect 5408 6808 5414 6820
rect 5445 6817 5457 6820
rect 5491 6817 5503 6851
rect 5445 6811 5503 6817
rect 5460 6780 5488 6811
rect 9766 6808 9772 6860
rect 9824 6848 9830 6860
rect 10045 6851 10103 6857
rect 10045 6848 10057 6851
rect 9824 6820 10057 6848
rect 9824 6808 9830 6820
rect 10045 6817 10057 6820
rect 10091 6817 10103 6851
rect 10045 6811 10103 6817
rect 10152 6820 13400 6848
rect 6914 6780 6920 6792
rect 5460 6752 6920 6780
rect 6914 6740 6920 6752
rect 6972 6740 6978 6792
rect 9582 6740 9588 6792
rect 9640 6780 9646 6792
rect 10152 6780 10180 6820
rect 9640 6752 10180 6780
rect 10505 6783 10563 6789
rect 9640 6740 9646 6752
rect 10505 6749 10517 6783
rect 10551 6749 10563 6783
rect 10505 6743 10563 6749
rect 5712 6715 5770 6721
rect 5712 6681 5724 6715
rect 5758 6712 5770 6715
rect 5810 6712 5816 6724
rect 5758 6684 5816 6712
rect 5758 6681 5770 6684
rect 5712 6675 5770 6681
rect 5810 6672 5816 6684
rect 5868 6672 5874 6724
rect 5902 6672 5908 6724
rect 5960 6712 5966 6724
rect 7162 6715 7220 6721
rect 7162 6712 7174 6715
rect 5960 6684 7174 6712
rect 5960 6672 5966 6684
rect 7162 6681 7174 6684
rect 7208 6681 7220 6715
rect 9953 6715 10011 6721
rect 9953 6712 9965 6715
rect 7162 6675 7220 6681
rect 9784 6684 9965 6712
rect 9784 6656 9812 6684
rect 9953 6681 9965 6684
rect 9999 6681 10011 6715
rect 9953 6675 10011 6681
rect 10042 6672 10048 6724
rect 10100 6712 10106 6724
rect 10520 6712 10548 6743
rect 10870 6740 10876 6792
rect 10928 6740 10934 6792
rect 13173 6783 13231 6789
rect 13173 6780 13185 6783
rect 12820 6752 13185 6780
rect 10100 6684 10548 6712
rect 10100 6672 10106 6684
rect 6638 6604 6644 6656
rect 6696 6644 6702 6656
rect 6825 6647 6883 6653
rect 6825 6644 6837 6647
rect 6696 6616 6837 6644
rect 6696 6604 6702 6616
rect 6825 6613 6837 6616
rect 6871 6613 6883 6647
rect 6825 6607 6883 6613
rect 8294 6604 8300 6656
rect 8352 6604 8358 6656
rect 9766 6604 9772 6656
rect 9824 6604 9830 6656
rect 9861 6647 9919 6653
rect 9861 6613 9873 6647
rect 9907 6644 9919 6647
rect 10888 6644 10916 6740
rect 12820 6724 12848 6752
rect 13173 6749 13185 6752
rect 13219 6749 13231 6783
rect 13173 6743 13231 6749
rect 13262 6740 13268 6792
rect 13320 6740 13326 6792
rect 13372 6780 13400 6820
rect 13446 6808 13452 6860
rect 13504 6848 13510 6860
rect 13504 6820 14136 6848
rect 13504 6808 13510 6820
rect 13538 6780 13544 6792
rect 13372 6752 13544 6780
rect 13538 6740 13544 6752
rect 13596 6740 13602 6792
rect 14108 6789 14136 6820
rect 16666 6808 16672 6860
rect 16724 6808 16730 6860
rect 14093 6783 14151 6789
rect 14093 6749 14105 6783
rect 14139 6780 14151 6783
rect 16684 6780 16712 6808
rect 17144 6789 17172 6888
rect 19426 6876 19432 6928
rect 19484 6916 19490 6928
rect 21726 6916 21732 6928
rect 19484 6888 21732 6916
rect 19484 6876 19490 6888
rect 21726 6876 21732 6888
rect 21784 6916 21790 6928
rect 22186 6916 22192 6928
rect 21784 6888 22192 6916
rect 21784 6876 21790 6888
rect 22186 6876 22192 6888
rect 22244 6916 22250 6928
rect 22244 6888 26372 6916
rect 22244 6876 22250 6888
rect 20806 6808 20812 6860
rect 20864 6848 20870 6860
rect 24949 6851 25007 6857
rect 24949 6848 24961 6851
rect 20864 6820 24961 6848
rect 20864 6808 20870 6820
rect 24949 6817 24961 6820
rect 24995 6817 25007 6851
rect 24949 6811 25007 6817
rect 14139 6752 16712 6780
rect 17129 6783 17187 6789
rect 14139 6749 14151 6752
rect 14093 6743 14151 6749
rect 17129 6749 17141 6783
rect 17175 6780 17187 6783
rect 17678 6780 17684 6792
rect 17175 6752 17684 6780
rect 17175 6749 17187 6752
rect 17129 6743 17187 6749
rect 17678 6740 17684 6752
rect 17736 6740 17742 6792
rect 19150 6740 19156 6792
rect 19208 6780 19214 6792
rect 23937 6783 23995 6789
rect 19208 6752 22048 6780
rect 19208 6740 19214 6752
rect 12802 6672 12808 6724
rect 12860 6672 12866 6724
rect 13280 6712 13308 6740
rect 22020 6724 22048 6752
rect 23937 6749 23949 6783
rect 23983 6780 23995 6783
rect 24118 6780 24124 6792
rect 23983 6752 24124 6780
rect 23983 6749 23995 6752
rect 23937 6743 23995 6749
rect 24118 6740 24124 6752
rect 24176 6740 24182 6792
rect 24228 6752 25360 6780
rect 13357 6715 13415 6721
rect 13357 6712 13369 6715
rect 13280 6684 13369 6712
rect 13357 6681 13369 6684
rect 13403 6681 13415 6715
rect 13357 6675 13415 6681
rect 13449 6715 13507 6721
rect 13449 6681 13461 6715
rect 13495 6712 13507 6715
rect 13906 6712 13912 6724
rect 13495 6684 13912 6712
rect 13495 6681 13507 6684
rect 13449 6675 13507 6681
rect 13906 6672 13912 6684
rect 13964 6672 13970 6724
rect 13998 6672 14004 6724
rect 14056 6712 14062 6724
rect 14338 6715 14396 6721
rect 14338 6712 14350 6715
rect 14056 6684 14350 6712
rect 14056 6672 14062 6684
rect 14338 6681 14350 6684
rect 14384 6681 14396 6715
rect 14338 6675 14396 6681
rect 16669 6715 16727 6721
rect 16669 6681 16681 6715
rect 16715 6712 16727 6715
rect 20622 6712 20628 6724
rect 16715 6684 20628 6712
rect 16715 6681 16727 6684
rect 16669 6675 16727 6681
rect 9907 6616 10916 6644
rect 9907 6613 9919 6616
rect 9861 6607 9919 6613
rect 12158 6604 12164 6656
rect 12216 6644 12222 6656
rect 16684 6644 16712 6675
rect 20622 6672 20628 6684
rect 20680 6672 20686 6724
rect 22002 6672 22008 6724
rect 22060 6712 22066 6724
rect 24228 6712 24256 6752
rect 22060 6684 24256 6712
rect 22060 6672 22066 6684
rect 24670 6672 24676 6724
rect 24728 6672 24734 6724
rect 24765 6715 24823 6721
rect 24765 6681 24777 6715
rect 24811 6712 24823 6715
rect 25225 6715 25283 6721
rect 25225 6712 25237 6715
rect 24811 6684 25237 6712
rect 24811 6681 24823 6684
rect 24765 6675 24823 6681
rect 25225 6681 25237 6684
rect 25271 6681 25283 6715
rect 25332 6712 25360 6752
rect 25498 6740 25504 6792
rect 25556 6780 25562 6792
rect 26344 6789 26372 6888
rect 25777 6783 25835 6789
rect 25777 6780 25789 6783
rect 25556 6752 25789 6780
rect 25556 6740 25562 6752
rect 25777 6749 25789 6752
rect 25823 6780 25835 6783
rect 25961 6783 26019 6789
rect 25961 6780 25973 6783
rect 25823 6752 25973 6780
rect 25823 6749 25835 6752
rect 25777 6743 25835 6749
rect 25961 6749 25973 6752
rect 26007 6749 26019 6783
rect 25961 6743 26019 6749
rect 26329 6783 26387 6789
rect 26329 6749 26341 6783
rect 26375 6749 26387 6783
rect 26329 6743 26387 6749
rect 26145 6715 26203 6721
rect 26145 6712 26157 6715
rect 25332 6684 26157 6712
rect 25225 6675 25283 6681
rect 26145 6681 26157 6684
rect 26191 6681 26203 6715
rect 26145 6675 26203 6681
rect 26237 6715 26295 6721
rect 26237 6681 26249 6715
rect 26283 6681 26295 6715
rect 26237 6675 26295 6681
rect 12216 6616 16712 6644
rect 12216 6604 12222 6616
rect 16758 6604 16764 6656
rect 16816 6604 16822 6656
rect 17310 6604 17316 6656
rect 17368 6644 17374 6656
rect 18782 6644 18788 6656
rect 17368 6616 18788 6644
rect 17368 6604 17374 6616
rect 18782 6604 18788 6616
rect 18840 6604 18846 6656
rect 19058 6604 19064 6656
rect 19116 6644 19122 6656
rect 21818 6644 21824 6656
rect 19116 6616 21824 6644
rect 19116 6604 19122 6616
rect 21818 6604 21824 6616
rect 21876 6604 21882 6656
rect 24026 6604 24032 6656
rect 24084 6644 24090 6656
rect 24121 6647 24179 6653
rect 24121 6644 24133 6647
rect 24084 6616 24133 6644
rect 24084 6604 24090 6616
rect 24121 6613 24133 6616
rect 24167 6613 24179 6647
rect 24121 6607 24179 6613
rect 24210 6604 24216 6656
rect 24268 6644 24274 6656
rect 24397 6647 24455 6653
rect 24397 6644 24409 6647
rect 24268 6616 24409 6644
rect 24268 6604 24274 6616
rect 24397 6613 24409 6616
rect 24443 6613 24455 6647
rect 24688 6644 24716 6672
rect 24857 6647 24915 6653
rect 24857 6644 24869 6647
rect 24688 6616 24869 6644
rect 24397 6607 24455 6613
rect 24857 6613 24869 6616
rect 24903 6613 24915 6647
rect 24857 6607 24915 6613
rect 25774 6604 25780 6656
rect 25832 6644 25838 6656
rect 26252 6644 26280 6675
rect 25832 6616 26280 6644
rect 25832 6604 25838 6616
rect 26418 6604 26424 6656
rect 26476 6644 26482 6656
rect 26513 6647 26571 6653
rect 26513 6644 26525 6647
rect 26476 6616 26525 6644
rect 26476 6604 26482 6616
rect 26513 6613 26525 6616
rect 26559 6613 26571 6647
rect 26513 6607 26571 6613
rect 1104 6554 31832 6576
rect 1104 6502 4922 6554
rect 4974 6502 4986 6554
rect 5038 6502 5050 6554
rect 5102 6502 5114 6554
rect 5166 6502 5178 6554
rect 5230 6502 5242 6554
rect 5294 6502 10922 6554
rect 10974 6502 10986 6554
rect 11038 6502 11050 6554
rect 11102 6502 11114 6554
rect 11166 6502 11178 6554
rect 11230 6502 11242 6554
rect 11294 6502 16922 6554
rect 16974 6502 16986 6554
rect 17038 6502 17050 6554
rect 17102 6502 17114 6554
rect 17166 6502 17178 6554
rect 17230 6502 17242 6554
rect 17294 6502 22922 6554
rect 22974 6502 22986 6554
rect 23038 6502 23050 6554
rect 23102 6502 23114 6554
rect 23166 6502 23178 6554
rect 23230 6502 23242 6554
rect 23294 6502 28922 6554
rect 28974 6502 28986 6554
rect 29038 6502 29050 6554
rect 29102 6502 29114 6554
rect 29166 6502 29178 6554
rect 29230 6502 29242 6554
rect 29294 6502 31832 6554
rect 1104 6480 31832 6502
rect 1581 6443 1639 6449
rect 1581 6409 1593 6443
rect 1627 6440 1639 6443
rect 4614 6440 4620 6452
rect 1627 6412 4620 6440
rect 1627 6409 1639 6412
rect 1581 6403 1639 6409
rect 4614 6400 4620 6412
rect 4672 6440 4678 6452
rect 5350 6440 5356 6452
rect 4672 6412 5356 6440
rect 4672 6400 4678 6412
rect 5350 6400 5356 6412
rect 5408 6400 5414 6452
rect 5902 6400 5908 6452
rect 5960 6400 5966 6452
rect 6181 6443 6239 6449
rect 6181 6409 6193 6443
rect 6227 6409 6239 6443
rect 6181 6403 6239 6409
rect 6196 6372 6224 6403
rect 7190 6400 7196 6452
rect 7248 6400 7254 6452
rect 7745 6443 7803 6449
rect 7745 6409 7757 6443
rect 7791 6440 7803 6443
rect 9125 6443 9183 6449
rect 7791 6412 8616 6440
rect 7791 6409 7803 6412
rect 7745 6403 7803 6409
rect 6610 6375 6668 6381
rect 6610 6372 6622 6375
rect 6196 6344 6622 6372
rect 6610 6341 6622 6344
rect 6656 6341 6668 6375
rect 6610 6335 6668 6341
rect 934 6264 940 6316
rect 992 6304 998 6316
rect 1397 6307 1455 6313
rect 1397 6304 1409 6307
rect 992 6276 1409 6304
rect 992 6264 998 6276
rect 1397 6273 1409 6276
rect 1443 6273 1455 6307
rect 1397 6267 1455 6273
rect 5442 6264 5448 6316
rect 5500 6264 5506 6316
rect 5718 6264 5724 6316
rect 5776 6264 5782 6316
rect 5997 6307 6055 6313
rect 5997 6273 6009 6307
rect 6043 6304 6055 6307
rect 7208 6304 7236 6400
rect 8588 6316 8616 6412
rect 9125 6409 9137 6443
rect 9171 6440 9183 6443
rect 9214 6440 9220 6452
rect 9171 6412 9220 6440
rect 9171 6409 9183 6412
rect 9125 6403 9183 6409
rect 9214 6400 9220 6412
rect 9272 6400 9278 6452
rect 11977 6443 12035 6449
rect 11977 6409 11989 6443
rect 12023 6409 12035 6443
rect 11977 6403 12035 6409
rect 6043 6276 7236 6304
rect 6043 6273 6055 6276
rect 5997 6267 6055 6273
rect 8294 6264 8300 6316
rect 8352 6304 8358 6316
rect 8389 6307 8447 6313
rect 8389 6304 8401 6307
rect 8352 6276 8401 6304
rect 8352 6264 8358 6276
rect 8389 6273 8401 6276
rect 8435 6273 8447 6307
rect 8389 6267 8447 6273
rect 8570 6264 8576 6316
rect 8628 6264 8634 6316
rect 8757 6307 8815 6313
rect 8757 6273 8769 6307
rect 8803 6273 8815 6307
rect 8757 6267 8815 6273
rect 5460 6236 5488 6264
rect 6365 6239 6423 6245
rect 6365 6236 6377 6239
rect 5460 6208 6377 6236
rect 6365 6205 6377 6208
rect 6411 6205 6423 6239
rect 6365 6199 6423 6205
rect 8478 6196 8484 6248
rect 8536 6236 8542 6248
rect 8772 6236 8800 6267
rect 8846 6264 8852 6316
rect 8904 6264 8910 6316
rect 8938 6264 8944 6316
rect 8996 6304 9002 6316
rect 9582 6304 9588 6316
rect 8996 6276 9588 6304
rect 8996 6264 9002 6276
rect 9582 6264 9588 6276
rect 9640 6264 9646 6316
rect 11885 6307 11943 6313
rect 11885 6273 11897 6307
rect 11931 6304 11943 6307
rect 11992 6304 12020 6403
rect 12250 6400 12256 6452
rect 12308 6440 12314 6452
rect 12437 6443 12495 6449
rect 12437 6440 12449 6443
rect 12308 6412 12449 6440
rect 12308 6400 12314 6412
rect 12437 6409 12449 6412
rect 12483 6409 12495 6443
rect 12437 6403 12495 6409
rect 12526 6400 12532 6452
rect 12584 6440 12590 6452
rect 12584 6412 13769 6440
rect 12584 6400 12590 6412
rect 13262 6372 13268 6384
rect 11931 6276 12020 6304
rect 12084 6344 13268 6372
rect 11931 6273 11943 6276
rect 11885 6267 11943 6273
rect 12084 6236 12112 6344
rect 13262 6332 13268 6344
rect 13320 6332 13326 6384
rect 12158 6264 12164 6316
rect 12216 6264 12222 6316
rect 12345 6307 12403 6313
rect 12345 6273 12357 6307
rect 12391 6304 12403 6307
rect 12805 6307 12863 6313
rect 12805 6304 12817 6307
rect 12391 6276 12817 6304
rect 12391 6273 12403 6276
rect 12345 6267 12403 6273
rect 12805 6273 12817 6276
rect 12851 6273 12863 6307
rect 12805 6267 12863 6273
rect 8536 6208 12112 6236
rect 8536 6196 8542 6208
rect 7466 6128 7472 6180
rect 7524 6168 7530 6180
rect 12176 6168 12204 6264
rect 12529 6239 12587 6245
rect 12529 6205 12541 6239
rect 12575 6205 12587 6239
rect 13357 6239 13415 6245
rect 13357 6236 13369 6239
rect 12529 6199 12587 6205
rect 12820 6208 13369 6236
rect 12544 6168 12572 6199
rect 7524 6140 12204 6168
rect 12406 6140 12572 6168
rect 7524 6128 7530 6140
rect 7834 6060 7840 6112
rect 7892 6060 7898 6112
rect 11698 6060 11704 6112
rect 11756 6060 11762 6112
rect 12066 6060 12072 6112
rect 12124 6100 12130 6112
rect 12406 6100 12434 6140
rect 12820 6112 12848 6208
rect 13357 6205 13369 6208
rect 13403 6205 13415 6239
rect 13741 6236 13769 6412
rect 13998 6400 14004 6452
rect 14056 6400 14062 6452
rect 14642 6400 14648 6452
rect 14700 6400 14706 6452
rect 17678 6400 17684 6452
rect 17736 6400 17742 6452
rect 19150 6400 19156 6452
rect 19208 6400 19214 6452
rect 19518 6400 19524 6452
rect 19576 6400 19582 6452
rect 19702 6400 19708 6452
rect 19760 6440 19766 6452
rect 22373 6443 22431 6449
rect 19760 6412 22324 6440
rect 19760 6400 19766 6412
rect 13817 6307 13875 6313
rect 13817 6273 13829 6307
rect 13863 6304 13875 6307
rect 14660 6304 14688 6400
rect 19058 6372 19064 6384
rect 13863 6276 14688 6304
rect 16776 6344 19064 6372
rect 13863 6273 13875 6276
rect 13817 6267 13875 6273
rect 16776 6248 16804 6344
rect 19058 6332 19064 6344
rect 19116 6332 19122 6384
rect 19168 6313 19196 6400
rect 19242 6381 19248 6384
rect 19241 6335 19248 6381
rect 19300 6372 19306 6384
rect 19300 6344 19341 6372
rect 19242 6332 19248 6335
rect 19300 6332 19306 6344
rect 22002 6332 22008 6384
rect 22060 6332 22066 6384
rect 17589 6307 17647 6313
rect 17589 6273 17601 6307
rect 17635 6304 17647 6307
rect 18049 6307 18107 6313
rect 18049 6304 18061 6307
rect 17635 6276 18061 6304
rect 17635 6273 17647 6276
rect 17589 6267 17647 6273
rect 18049 6273 18061 6276
rect 18095 6273 18107 6307
rect 18969 6307 19027 6313
rect 18969 6304 18981 6307
rect 18049 6267 18107 6273
rect 18616 6276 18981 6304
rect 16758 6236 16764 6248
rect 13741 6208 16764 6236
rect 13357 6199 13415 6205
rect 16758 6196 16764 6208
rect 16816 6196 16822 6248
rect 17862 6196 17868 6248
rect 17920 6196 17926 6248
rect 18616 6245 18644 6276
rect 18969 6273 18981 6276
rect 19015 6273 19027 6307
rect 18969 6267 19027 6273
rect 19153 6307 19211 6313
rect 19153 6273 19165 6307
rect 19199 6273 19211 6307
rect 19153 6267 19211 6273
rect 19380 6264 19386 6316
rect 19438 6264 19444 6316
rect 21821 6307 21879 6313
rect 21821 6304 21833 6307
rect 21560 6276 21833 6304
rect 21560 6248 21588 6276
rect 21821 6273 21833 6276
rect 21867 6273 21879 6307
rect 21821 6267 21879 6273
rect 22094 6264 22100 6316
rect 22152 6264 22158 6316
rect 22186 6264 22192 6316
rect 22244 6264 22250 6316
rect 22296 6304 22324 6412
rect 22373 6409 22385 6443
rect 22419 6440 22431 6443
rect 22646 6440 22652 6452
rect 22419 6412 22652 6440
rect 22419 6409 22431 6412
rect 22373 6403 22431 6409
rect 22646 6400 22652 6412
rect 22704 6400 22710 6452
rect 23750 6400 23756 6452
rect 23808 6440 23814 6452
rect 23808 6412 23960 6440
rect 23808 6400 23814 6412
rect 23932 6381 23960 6412
rect 24118 6400 24124 6452
rect 24176 6440 24182 6452
rect 25133 6443 25191 6449
rect 25133 6440 25145 6443
rect 24176 6412 25145 6440
rect 24176 6400 24182 6412
rect 25133 6409 25145 6412
rect 25179 6409 25191 6443
rect 25133 6403 25191 6409
rect 23928 6375 23986 6381
rect 23928 6341 23940 6375
rect 23974 6341 23986 6375
rect 25590 6372 25596 6384
rect 23928 6335 23986 6341
rect 25424 6344 25596 6372
rect 25424 6304 25452 6344
rect 25590 6332 25596 6344
rect 25648 6332 25654 6384
rect 22296 6276 25452 6304
rect 25501 6307 25559 6313
rect 25501 6273 25513 6307
rect 25547 6304 25559 6307
rect 25961 6307 26019 6313
rect 25961 6304 25973 6307
rect 25547 6276 25973 6304
rect 25547 6273 25559 6276
rect 25501 6267 25559 6273
rect 25961 6273 25973 6276
rect 26007 6273 26019 6307
rect 25961 6267 26019 6273
rect 18601 6239 18659 6245
rect 18601 6236 18613 6239
rect 18248 6208 18613 6236
rect 18248 6112 18276 6208
rect 18601 6205 18613 6208
rect 18647 6205 18659 6239
rect 18601 6199 18659 6205
rect 21542 6196 21548 6248
rect 21600 6196 21606 6248
rect 23658 6196 23664 6248
rect 23716 6196 23722 6248
rect 25685 6239 25743 6245
rect 25685 6205 25697 6239
rect 25731 6205 25743 6239
rect 26513 6239 26571 6245
rect 26513 6236 26525 6239
rect 25685 6199 25743 6205
rect 25792 6208 26525 6236
rect 25041 6171 25099 6177
rect 25041 6137 25053 6171
rect 25087 6168 25099 6171
rect 25498 6168 25504 6180
rect 25087 6140 25504 6168
rect 25087 6137 25099 6140
rect 25041 6131 25099 6137
rect 25498 6128 25504 6140
rect 25556 6128 25562 6180
rect 12124 6072 12434 6100
rect 12124 6060 12130 6072
rect 12802 6060 12808 6112
rect 12860 6060 12866 6112
rect 17221 6103 17279 6109
rect 17221 6069 17233 6103
rect 17267 6100 17279 6103
rect 17402 6100 17408 6112
rect 17267 6072 17408 6100
rect 17267 6069 17279 6072
rect 17221 6063 17279 6069
rect 17402 6060 17408 6072
rect 17460 6060 17466 6112
rect 18230 6060 18236 6112
rect 18288 6060 18294 6112
rect 20990 6060 20996 6112
rect 21048 6060 21054 6112
rect 23566 6060 23572 6112
rect 23624 6100 23630 6112
rect 25700 6100 25728 6199
rect 25792 6112 25820 6208
rect 26513 6205 26525 6208
rect 26559 6205 26571 6239
rect 26513 6199 26571 6205
rect 23624 6072 25728 6100
rect 23624 6060 23630 6072
rect 25774 6060 25780 6112
rect 25832 6060 25838 6112
rect 1104 6010 31832 6032
rect 1104 5958 4182 6010
rect 4234 5958 4246 6010
rect 4298 5958 4310 6010
rect 4362 5958 4374 6010
rect 4426 5958 4438 6010
rect 4490 5958 4502 6010
rect 4554 5958 10182 6010
rect 10234 5958 10246 6010
rect 10298 5958 10310 6010
rect 10362 5958 10374 6010
rect 10426 5958 10438 6010
rect 10490 5958 10502 6010
rect 10554 5958 16182 6010
rect 16234 5958 16246 6010
rect 16298 5958 16310 6010
rect 16362 5958 16374 6010
rect 16426 5958 16438 6010
rect 16490 5958 16502 6010
rect 16554 5958 22182 6010
rect 22234 5958 22246 6010
rect 22298 5958 22310 6010
rect 22362 5958 22374 6010
rect 22426 5958 22438 6010
rect 22490 5958 22502 6010
rect 22554 5958 28182 6010
rect 28234 5958 28246 6010
rect 28298 5958 28310 6010
rect 28362 5958 28374 6010
rect 28426 5958 28438 6010
rect 28490 5958 28502 6010
rect 28554 5958 31832 6010
rect 1104 5936 31832 5958
rect 5718 5856 5724 5908
rect 5776 5896 5782 5908
rect 6181 5899 6239 5905
rect 6181 5896 6193 5899
rect 5776 5868 6193 5896
rect 5776 5856 5782 5868
rect 6181 5865 6193 5868
rect 6227 5865 6239 5899
rect 6181 5859 6239 5865
rect 7834 5856 7840 5908
rect 7892 5856 7898 5908
rect 11606 5896 11612 5908
rect 11440 5868 11612 5896
rect 6825 5763 6883 5769
rect 6825 5729 6837 5763
rect 6871 5760 6883 5763
rect 7742 5760 7748 5772
rect 6871 5732 7748 5760
rect 6871 5729 6883 5732
rect 6825 5723 6883 5729
rect 7742 5720 7748 5732
rect 7800 5720 7806 5772
rect 6549 5695 6607 5701
rect 6549 5661 6561 5695
rect 6595 5692 6607 5695
rect 7852 5692 7880 5856
rect 11440 5769 11468 5868
rect 11606 5856 11612 5868
rect 11664 5856 11670 5908
rect 12802 5856 12808 5908
rect 12860 5856 12866 5908
rect 18230 5856 18236 5908
rect 18288 5856 18294 5908
rect 18892 5868 20852 5896
rect 18892 5828 18920 5868
rect 17880 5800 18920 5828
rect 18984 5800 20484 5828
rect 17880 5772 17908 5800
rect 11425 5763 11483 5769
rect 11425 5729 11437 5763
rect 11471 5729 11483 5763
rect 11425 5723 11483 5729
rect 6595 5664 7880 5692
rect 11440 5692 11468 5723
rect 13906 5720 13912 5772
rect 13964 5720 13970 5772
rect 14274 5720 14280 5772
rect 14332 5760 14338 5772
rect 14645 5763 14703 5769
rect 14645 5760 14657 5763
rect 14332 5732 14657 5760
rect 14332 5720 14338 5732
rect 14645 5729 14657 5732
rect 14691 5729 14703 5763
rect 14645 5723 14703 5729
rect 16666 5720 16672 5772
rect 16724 5760 16730 5772
rect 16853 5763 16911 5769
rect 16853 5760 16865 5763
rect 16724 5732 16865 5760
rect 16724 5720 16730 5732
rect 16853 5729 16865 5732
rect 16899 5729 16911 5763
rect 16853 5723 16911 5729
rect 17862 5720 17868 5772
rect 17920 5720 17926 5772
rect 18782 5720 18788 5772
rect 18840 5720 18846 5772
rect 18984 5769 19012 5800
rect 18969 5763 19027 5769
rect 18969 5729 18981 5763
rect 19015 5729 19027 5763
rect 18969 5723 19027 5729
rect 19242 5720 19248 5772
rect 19300 5720 19306 5772
rect 12158 5692 12164 5704
rect 11440 5664 12164 5692
rect 6595 5661 6607 5664
rect 6549 5655 6607 5661
rect 12158 5652 12164 5664
rect 12216 5692 12222 5704
rect 12802 5692 12808 5704
rect 12216 5664 12808 5692
rect 12216 5652 12222 5664
rect 12802 5652 12808 5664
rect 12860 5652 12866 5704
rect 13924 5692 13952 5720
rect 15473 5695 15531 5701
rect 15473 5692 15485 5695
rect 13924 5664 15485 5692
rect 15473 5661 15485 5664
rect 15519 5661 15531 5695
rect 15473 5655 15531 5661
rect 18874 5652 18880 5704
rect 18932 5692 18938 5704
rect 19260 5692 19288 5720
rect 19889 5695 19947 5701
rect 19889 5692 19901 5695
rect 18932 5664 19901 5692
rect 18932 5652 18938 5664
rect 19889 5661 19901 5664
rect 19935 5661 19947 5695
rect 19889 5655 19947 5661
rect 5350 5584 5356 5636
rect 5408 5624 5414 5636
rect 6641 5627 6699 5633
rect 6641 5624 6653 5627
rect 5408 5596 6653 5624
rect 5408 5584 5414 5596
rect 6641 5593 6653 5596
rect 6687 5624 6699 5627
rect 7466 5624 7472 5636
rect 6687 5596 7472 5624
rect 6687 5593 6699 5596
rect 6641 5587 6699 5593
rect 7466 5584 7472 5596
rect 7524 5584 7530 5636
rect 11698 5633 11704 5636
rect 11692 5624 11704 5633
rect 11659 5596 11704 5624
rect 11692 5587 11704 5596
rect 11698 5584 11704 5587
rect 11756 5584 11762 5636
rect 14461 5627 14519 5633
rect 14461 5593 14473 5627
rect 14507 5624 14519 5627
rect 14921 5627 14979 5633
rect 14921 5624 14933 5627
rect 14507 5596 14933 5624
rect 14507 5593 14519 5596
rect 14461 5587 14519 5593
rect 14921 5593 14933 5596
rect 14967 5593 14979 5627
rect 14921 5587 14979 5593
rect 17120 5627 17178 5633
rect 17120 5593 17132 5627
rect 17166 5624 17178 5627
rect 17310 5624 17316 5636
rect 17166 5596 17316 5624
rect 17166 5593 17178 5596
rect 17120 5587 17178 5593
rect 17310 5584 17316 5596
rect 17368 5584 17374 5636
rect 18693 5627 18751 5633
rect 17420 5596 18460 5624
rect 14090 5516 14096 5568
rect 14148 5516 14154 5568
rect 14553 5559 14611 5565
rect 14553 5525 14565 5559
rect 14599 5556 14611 5559
rect 15102 5556 15108 5568
rect 14599 5528 15108 5556
rect 14599 5525 14611 5528
rect 14553 5519 14611 5525
rect 15102 5516 15108 5528
rect 15160 5556 15166 5568
rect 17420 5556 17448 5596
rect 15160 5528 17448 5556
rect 15160 5516 15166 5528
rect 18322 5516 18328 5568
rect 18380 5516 18386 5568
rect 18432 5556 18460 5596
rect 18693 5593 18705 5627
rect 18739 5624 18751 5627
rect 19245 5627 19303 5633
rect 19245 5624 19257 5627
rect 18739 5596 19257 5624
rect 18739 5593 18751 5596
rect 18693 5587 18751 5593
rect 19245 5593 19257 5596
rect 19291 5593 19303 5627
rect 20456 5624 20484 5800
rect 20824 5772 20852 5868
rect 20990 5856 20996 5908
rect 21048 5856 21054 5908
rect 21818 5856 21824 5908
rect 21876 5856 21882 5908
rect 23566 5856 23572 5908
rect 23624 5856 23630 5908
rect 23750 5856 23756 5908
rect 23808 5896 23814 5908
rect 23937 5899 23995 5905
rect 23937 5896 23949 5899
rect 23808 5868 23949 5896
rect 23808 5856 23814 5868
rect 23937 5865 23949 5868
rect 23983 5865 23995 5899
rect 23937 5859 23995 5865
rect 20622 5720 20628 5772
rect 20680 5720 20686 5772
rect 20806 5720 20812 5772
rect 20864 5720 20870 5772
rect 20533 5695 20591 5701
rect 20533 5661 20545 5695
rect 20579 5692 20591 5695
rect 21008 5692 21036 5856
rect 21634 5760 21640 5772
rect 20579 5664 21036 5692
rect 21100 5732 21640 5760
rect 20579 5661 20591 5664
rect 20533 5655 20591 5661
rect 21100 5624 21128 5732
rect 21634 5720 21640 5732
rect 21692 5720 21698 5772
rect 21729 5763 21787 5769
rect 21729 5729 21741 5763
rect 21775 5760 21787 5763
rect 21836 5760 21864 5856
rect 21775 5732 21864 5760
rect 21775 5729 21787 5732
rect 21729 5723 21787 5729
rect 21910 5720 21916 5772
rect 21968 5760 21974 5772
rect 23584 5760 23612 5856
rect 25774 5788 25780 5840
rect 25832 5788 25838 5840
rect 21968 5732 23612 5760
rect 21968 5720 21974 5732
rect 23658 5720 23664 5772
rect 23716 5760 23722 5772
rect 24397 5763 24455 5769
rect 24397 5760 24409 5763
rect 23716 5732 24409 5760
rect 23716 5720 23722 5732
rect 24397 5729 24409 5732
rect 24443 5729 24455 5763
rect 24397 5723 24455 5729
rect 24026 5652 24032 5704
rect 24084 5652 24090 5704
rect 24121 5695 24179 5701
rect 24121 5661 24133 5695
rect 24167 5692 24179 5695
rect 24210 5692 24216 5704
rect 24167 5664 24216 5692
rect 24167 5661 24179 5664
rect 24121 5655 24179 5661
rect 24210 5652 24216 5664
rect 24268 5652 24274 5704
rect 20456 5596 21128 5624
rect 24044 5624 24072 5652
rect 24642 5627 24700 5633
rect 24642 5624 24654 5627
rect 24044 5596 24654 5624
rect 19245 5587 19303 5593
rect 24642 5593 24654 5596
rect 24688 5593 24700 5627
rect 24642 5587 24700 5593
rect 19702 5556 19708 5568
rect 18432 5528 19708 5556
rect 19702 5516 19708 5528
rect 19760 5516 19766 5568
rect 19794 5516 19800 5568
rect 19852 5556 19858 5568
rect 20165 5559 20223 5565
rect 20165 5556 20177 5559
rect 19852 5528 20177 5556
rect 19852 5516 19858 5528
rect 20165 5525 20177 5528
rect 20211 5525 20223 5559
rect 20165 5519 20223 5525
rect 21266 5516 21272 5568
rect 21324 5516 21330 5568
rect 21634 5516 21640 5568
rect 21692 5516 21698 5568
rect 1104 5466 31832 5488
rect 1104 5414 4922 5466
rect 4974 5414 4986 5466
rect 5038 5414 5050 5466
rect 5102 5414 5114 5466
rect 5166 5414 5178 5466
rect 5230 5414 5242 5466
rect 5294 5414 10922 5466
rect 10974 5414 10986 5466
rect 11038 5414 11050 5466
rect 11102 5414 11114 5466
rect 11166 5414 11178 5466
rect 11230 5414 11242 5466
rect 11294 5414 16922 5466
rect 16974 5414 16986 5466
rect 17038 5414 17050 5466
rect 17102 5414 17114 5466
rect 17166 5414 17178 5466
rect 17230 5414 17242 5466
rect 17294 5414 22922 5466
rect 22974 5414 22986 5466
rect 23038 5414 23050 5466
rect 23102 5414 23114 5466
rect 23166 5414 23178 5466
rect 23230 5414 23242 5466
rect 23294 5414 28922 5466
rect 28974 5414 28986 5466
rect 29038 5414 29050 5466
rect 29102 5414 29114 5466
rect 29166 5414 29178 5466
rect 29230 5414 29242 5466
rect 29294 5414 31832 5466
rect 1104 5392 31832 5414
rect 8113 5355 8171 5361
rect 8113 5321 8125 5355
rect 8159 5352 8171 5355
rect 8662 5352 8668 5364
rect 8159 5324 8668 5352
rect 8159 5321 8171 5324
rect 8113 5315 8171 5321
rect 8662 5312 8668 5324
rect 8720 5312 8726 5364
rect 8757 5355 8815 5361
rect 8757 5321 8769 5355
rect 8803 5352 8815 5355
rect 9766 5352 9772 5364
rect 8803 5324 9772 5352
rect 8803 5321 8815 5324
rect 8757 5315 8815 5321
rect 9766 5312 9772 5324
rect 9824 5312 9830 5364
rect 13906 5312 13912 5364
rect 13964 5352 13970 5364
rect 14185 5355 14243 5361
rect 14185 5352 14197 5355
rect 13964 5324 14197 5352
rect 13964 5312 13970 5324
rect 14185 5321 14197 5324
rect 14231 5321 14243 5355
rect 14185 5315 14243 5321
rect 17129 5355 17187 5361
rect 17129 5321 17141 5355
rect 17175 5352 17187 5355
rect 17310 5352 17316 5364
rect 17175 5324 17316 5352
rect 17175 5321 17187 5324
rect 17129 5315 17187 5321
rect 17310 5312 17316 5324
rect 17368 5312 17374 5364
rect 17402 5312 17408 5364
rect 17460 5312 17466 5364
rect 18874 5312 18880 5364
rect 18932 5312 18938 5364
rect 19797 5355 19855 5361
rect 19797 5321 19809 5355
rect 19843 5352 19855 5355
rect 19843 5324 20024 5352
rect 19843 5321 19855 5324
rect 19797 5315 19855 5321
rect 14274 5284 14280 5296
rect 8680 5256 14280 5284
rect 8018 5176 8024 5228
rect 8076 5176 8082 5228
rect 8680 5157 8708 5256
rect 14274 5244 14280 5256
rect 14332 5244 14338 5296
rect 13078 5225 13084 5228
rect 8849 5219 8907 5225
rect 8849 5185 8861 5219
rect 8895 5216 8907 5219
rect 9309 5219 9367 5225
rect 9309 5216 9321 5219
rect 8895 5188 9321 5216
rect 8895 5185 8907 5188
rect 8849 5179 8907 5185
rect 9309 5185 9321 5188
rect 9355 5185 9367 5219
rect 9309 5179 9367 5185
rect 13072 5179 13084 5225
rect 13078 5176 13084 5179
rect 13136 5176 13142 5228
rect 17313 5219 17371 5225
rect 17313 5185 17325 5219
rect 17359 5216 17371 5219
rect 17420 5216 17448 5312
rect 19996 5284 20024 5324
rect 21266 5312 21272 5364
rect 21324 5312 21330 5364
rect 21634 5312 21640 5364
rect 21692 5352 21698 5364
rect 21913 5355 21971 5361
rect 21913 5352 21925 5355
rect 21692 5324 21925 5352
rect 21692 5312 21698 5324
rect 21913 5321 21925 5324
rect 21959 5321 21971 5355
rect 21913 5315 21971 5321
rect 20134 5287 20192 5293
rect 20134 5284 20146 5287
rect 17512 5256 19932 5284
rect 19996 5256 20146 5284
rect 17512 5225 17540 5256
rect 19904 5228 19932 5256
rect 20134 5253 20146 5256
rect 20180 5253 20192 5287
rect 20134 5247 20192 5253
rect 17770 5225 17776 5228
rect 17359 5188 17448 5216
rect 17497 5219 17555 5225
rect 17359 5185 17371 5188
rect 17313 5179 17371 5185
rect 17497 5185 17509 5219
rect 17543 5185 17555 5219
rect 17497 5179 17555 5185
rect 17764 5179 17776 5225
rect 17770 5176 17776 5179
rect 17828 5176 17834 5228
rect 19613 5219 19671 5225
rect 19613 5185 19625 5219
rect 19659 5216 19671 5219
rect 19794 5216 19800 5228
rect 19659 5188 19800 5216
rect 19659 5185 19671 5188
rect 19613 5179 19671 5185
rect 19794 5176 19800 5188
rect 19852 5176 19858 5228
rect 19886 5176 19892 5228
rect 19944 5176 19950 5228
rect 21284 5216 21312 5312
rect 21545 5219 21603 5225
rect 21545 5216 21557 5219
rect 21284 5188 21557 5216
rect 21545 5185 21557 5188
rect 21591 5185 21603 5219
rect 21545 5179 21603 5185
rect 22094 5176 22100 5228
rect 22152 5216 22158 5228
rect 22465 5219 22523 5225
rect 22465 5216 22477 5219
rect 22152 5188 22477 5216
rect 22152 5176 22158 5188
rect 22465 5185 22477 5188
rect 22511 5185 22523 5219
rect 22465 5179 22523 5185
rect 8297 5151 8355 5157
rect 8297 5117 8309 5151
rect 8343 5148 8355 5151
rect 8665 5151 8723 5157
rect 8665 5148 8677 5151
rect 8343 5120 8677 5148
rect 8343 5117 8355 5120
rect 8297 5111 8355 5117
rect 8665 5117 8677 5120
rect 8711 5117 8723 5151
rect 9861 5151 9919 5157
rect 9861 5148 9873 5151
rect 8665 5111 8723 5117
rect 8864 5120 9873 5148
rect 8864 5092 8892 5120
rect 9861 5117 9873 5120
rect 9907 5117 9919 5151
rect 9861 5111 9919 5117
rect 12802 5108 12808 5160
rect 12860 5108 12866 5160
rect 8846 5040 8852 5092
rect 8904 5040 8910 5092
rect 7282 4972 7288 5024
rect 7340 5012 7346 5024
rect 7653 5015 7711 5021
rect 7653 5012 7665 5015
rect 7340 4984 7665 5012
rect 7340 4972 7346 4984
rect 7653 4981 7665 4984
rect 7699 4981 7711 5015
rect 7653 4975 7711 4981
rect 9214 4972 9220 5024
rect 9272 4972 9278 5024
rect 12820 5012 12848 5108
rect 21269 5083 21327 5089
rect 21269 5049 21281 5083
rect 21315 5080 21327 5083
rect 21542 5080 21548 5092
rect 21315 5052 21548 5080
rect 21315 5049 21327 5052
rect 21269 5043 21327 5049
rect 21542 5040 21548 5052
rect 21600 5040 21606 5092
rect 15470 5012 15476 5024
rect 12820 4984 15476 5012
rect 15470 4972 15476 4984
rect 15528 4972 15534 5024
rect 21358 4972 21364 5024
rect 21416 4972 21422 5024
rect 1104 4922 31832 4944
rect 1104 4870 4182 4922
rect 4234 4870 4246 4922
rect 4298 4870 4310 4922
rect 4362 4870 4374 4922
rect 4426 4870 4438 4922
rect 4490 4870 4502 4922
rect 4554 4870 10182 4922
rect 10234 4870 10246 4922
rect 10298 4870 10310 4922
rect 10362 4870 10374 4922
rect 10426 4870 10438 4922
rect 10490 4870 10502 4922
rect 10554 4870 16182 4922
rect 16234 4870 16246 4922
rect 16298 4870 16310 4922
rect 16362 4870 16374 4922
rect 16426 4870 16438 4922
rect 16490 4870 16502 4922
rect 16554 4870 22182 4922
rect 22234 4870 22246 4922
rect 22298 4870 22310 4922
rect 22362 4870 22374 4922
rect 22426 4870 22438 4922
rect 22490 4870 22502 4922
rect 22554 4870 28182 4922
rect 28234 4870 28246 4922
rect 28298 4870 28310 4922
rect 28362 4870 28374 4922
rect 28426 4870 28438 4922
rect 28490 4870 28502 4922
rect 28554 4870 31832 4922
rect 1104 4848 31832 4870
rect 8018 4768 8024 4820
rect 8076 4808 8082 4820
rect 8941 4811 8999 4817
rect 8941 4808 8953 4811
rect 8076 4780 8953 4808
rect 8076 4768 8082 4780
rect 8941 4777 8953 4780
rect 8987 4777 8999 4811
rect 8941 4771 8999 4777
rect 9214 4768 9220 4820
rect 9272 4768 9278 4820
rect 13078 4768 13084 4820
rect 13136 4808 13142 4820
rect 13173 4811 13231 4817
rect 13173 4808 13185 4811
rect 13136 4780 13185 4808
rect 13136 4768 13142 4780
rect 13173 4777 13185 4780
rect 13219 4777 13231 4811
rect 13173 4771 13231 4777
rect 14090 4768 14096 4820
rect 14148 4768 14154 4820
rect 17770 4768 17776 4820
rect 17828 4808 17834 4820
rect 17865 4811 17923 4817
rect 17865 4808 17877 4811
rect 17828 4780 17877 4808
rect 17828 4768 17834 4780
rect 17865 4777 17877 4780
rect 17911 4777 17923 4811
rect 17865 4771 17923 4777
rect 22094 4768 22100 4820
rect 22152 4768 22158 4820
rect 8757 4743 8815 4749
rect 8757 4709 8769 4743
rect 8803 4740 8815 4743
rect 8846 4740 8852 4752
rect 8803 4712 8852 4740
rect 8803 4709 8815 4712
rect 8757 4703 8815 4709
rect 8846 4700 8852 4712
rect 8904 4700 8910 4752
rect 6914 4632 6920 4684
rect 6972 4672 6978 4684
rect 7377 4675 7435 4681
rect 7377 4672 7389 4675
rect 6972 4644 7389 4672
rect 6972 4632 6978 4644
rect 7377 4641 7389 4644
rect 7423 4641 7435 4675
rect 7377 4635 7435 4641
rect 8386 4632 8392 4684
rect 8444 4632 8450 4684
rect 9232 4672 9260 4768
rect 14108 4672 14136 4768
rect 9232 4644 9904 4672
rect 7101 4607 7159 4613
rect 7101 4573 7113 4607
rect 7147 4604 7159 4607
rect 7282 4604 7288 4616
rect 7147 4576 7288 4604
rect 7147 4573 7159 4576
rect 7101 4567 7159 4573
rect 7282 4564 7288 4576
rect 7340 4564 7346 4616
rect 8404 4604 8432 4632
rect 9876 4613 9904 4644
rect 13372 4644 14136 4672
rect 9493 4607 9551 4613
rect 9493 4604 9505 4607
rect 8404 4576 9505 4604
rect 9493 4573 9505 4576
rect 9539 4573 9551 4607
rect 9493 4567 9551 4573
rect 9861 4607 9919 4613
rect 9861 4573 9873 4607
rect 9907 4573 9919 4607
rect 9861 4567 9919 4573
rect 10778 4564 10784 4616
rect 10836 4604 10842 4616
rect 13372 4613 13400 4644
rect 15194 4632 15200 4684
rect 15252 4672 15258 4684
rect 15565 4675 15623 4681
rect 15565 4672 15577 4675
rect 15252 4644 15577 4672
rect 15252 4632 15258 4644
rect 15565 4641 15577 4644
rect 15611 4641 15623 4675
rect 15565 4635 15623 4641
rect 19886 4632 19892 4684
rect 19944 4672 19950 4684
rect 20717 4675 20775 4681
rect 20717 4672 20729 4675
rect 19944 4644 20729 4672
rect 19944 4632 19950 4644
rect 20717 4641 20729 4644
rect 20763 4641 20775 4675
rect 20717 4635 20775 4641
rect 11057 4607 11115 4613
rect 11057 4604 11069 4607
rect 10836 4576 11069 4604
rect 10836 4564 10842 4576
rect 11057 4573 11069 4576
rect 11103 4573 11115 4607
rect 11057 4567 11115 4573
rect 13357 4607 13415 4613
rect 13357 4573 13369 4607
rect 13403 4573 13415 4607
rect 13357 4567 13415 4573
rect 15289 4607 15347 4613
rect 15289 4573 15301 4607
rect 15335 4573 15347 4607
rect 15289 4567 15347 4573
rect 18049 4607 18107 4613
rect 18049 4573 18061 4607
rect 18095 4604 18107 4607
rect 18322 4604 18328 4616
rect 18095 4576 18328 4604
rect 18095 4573 18107 4576
rect 18049 4567 18107 4573
rect 7644 4539 7702 4545
rect 7644 4505 7656 4539
rect 7690 4536 7702 4539
rect 15304 4536 15332 4567
rect 18322 4564 18328 4576
rect 18380 4564 18386 4616
rect 20984 4607 21042 4613
rect 20984 4573 20996 4607
rect 21030 4604 21042 4607
rect 21358 4604 21364 4616
rect 21030 4576 21364 4604
rect 21030 4573 21042 4576
rect 20984 4567 21042 4573
rect 21358 4564 21364 4576
rect 21416 4564 21422 4616
rect 15470 4536 15476 4548
rect 7690 4508 9720 4536
rect 15304 4508 15476 4536
rect 7690 4505 7702 4508
rect 7644 4499 7702 4505
rect 7282 4428 7288 4480
rect 7340 4428 7346 4480
rect 9692 4477 9720 4508
rect 15470 4496 15476 4508
rect 15528 4496 15534 4548
rect 16574 4496 16580 4548
rect 16632 4496 16638 4548
rect 22066 4508 31248 4536
rect 9677 4471 9735 4477
rect 9677 4437 9689 4471
rect 9723 4437 9735 4471
rect 9677 4431 9735 4437
rect 10502 4428 10508 4480
rect 10560 4428 10566 4480
rect 15010 4428 15016 4480
rect 15068 4468 15074 4480
rect 17037 4471 17095 4477
rect 17037 4468 17049 4471
rect 15068 4440 17049 4468
rect 15068 4428 15074 4440
rect 17037 4437 17049 4440
rect 17083 4468 17095 4471
rect 22066 4468 22094 4508
rect 31220 4480 31248 4508
rect 17083 4440 22094 4468
rect 17083 4437 17095 4440
rect 17037 4431 17095 4437
rect 31202 4428 31208 4480
rect 31260 4428 31266 4480
rect 1104 4378 31832 4400
rect 1104 4326 4922 4378
rect 4974 4326 4986 4378
rect 5038 4326 5050 4378
rect 5102 4326 5114 4378
rect 5166 4326 5178 4378
rect 5230 4326 5242 4378
rect 5294 4326 10922 4378
rect 10974 4326 10986 4378
rect 11038 4326 11050 4378
rect 11102 4326 11114 4378
rect 11166 4326 11178 4378
rect 11230 4326 11242 4378
rect 11294 4326 16922 4378
rect 16974 4326 16986 4378
rect 17038 4326 17050 4378
rect 17102 4326 17114 4378
rect 17166 4326 17178 4378
rect 17230 4326 17242 4378
rect 17294 4326 22922 4378
rect 22974 4326 22986 4378
rect 23038 4326 23050 4378
rect 23102 4326 23114 4378
rect 23166 4326 23178 4378
rect 23230 4326 23242 4378
rect 23294 4326 28922 4378
rect 28974 4326 28986 4378
rect 29038 4326 29050 4378
rect 29102 4326 29114 4378
rect 29166 4326 29178 4378
rect 29230 4326 29242 4378
rect 29294 4326 31832 4378
rect 1104 4304 31832 4326
rect 7282 4224 7288 4276
rect 7340 4264 7346 4276
rect 7340 4236 7420 4264
rect 7340 4224 7346 4236
rect 7392 4205 7420 4236
rect 8386 4224 8392 4276
rect 8444 4264 8450 4276
rect 8481 4267 8539 4273
rect 8481 4264 8493 4267
rect 8444 4236 8493 4264
rect 8444 4224 8450 4236
rect 8481 4233 8493 4236
rect 8527 4233 8539 4267
rect 8481 4227 8539 4233
rect 10045 4267 10103 4273
rect 10045 4233 10057 4267
rect 10091 4264 10103 4267
rect 10502 4264 10508 4276
rect 10091 4236 10508 4264
rect 10091 4233 10103 4236
rect 10045 4227 10103 4233
rect 10502 4224 10508 4236
rect 10560 4224 10566 4276
rect 15010 4224 15016 4276
rect 15068 4224 15074 4276
rect 7368 4199 7426 4205
rect 7368 4165 7380 4199
rect 7414 4165 7426 4199
rect 7368 4159 7426 4165
rect 10873 4199 10931 4205
rect 10873 4165 10885 4199
rect 10919 4196 10931 4199
rect 11517 4199 11575 4205
rect 11517 4196 11529 4199
rect 10919 4168 11529 4196
rect 10919 4165 10931 4168
rect 10873 4159 10931 4165
rect 11517 4165 11529 4168
rect 11563 4165 11575 4199
rect 11517 4159 11575 4165
rect 15841 4199 15899 4205
rect 15841 4165 15853 4199
rect 15887 4196 15899 4199
rect 17402 4196 17408 4208
rect 15887 4168 17408 4196
rect 15887 4165 15899 4168
rect 15841 4159 15899 4165
rect 17402 4156 17408 4168
rect 17460 4156 17466 4208
rect 6914 4088 6920 4140
rect 6972 4128 6978 4140
rect 7101 4131 7159 4137
rect 7101 4128 7113 4131
rect 6972 4100 7113 4128
rect 6972 4088 6978 4100
rect 7101 4097 7113 4100
rect 7147 4097 7159 4131
rect 7101 4091 7159 4097
rect 10137 4131 10195 4137
rect 10137 4097 10149 4131
rect 10183 4128 10195 4131
rect 10183 4100 10548 4128
rect 10183 4097 10195 4100
rect 10137 4091 10195 4097
rect 10042 4020 10048 4072
rect 10100 4060 10106 4072
rect 10229 4063 10287 4069
rect 10229 4060 10241 4063
rect 10100 4032 10241 4060
rect 10100 4020 10106 4032
rect 10229 4029 10241 4032
rect 10275 4029 10287 4063
rect 10520 4060 10548 4100
rect 10594 4088 10600 4140
rect 10652 4128 10658 4140
rect 10965 4131 11023 4137
rect 10965 4128 10977 4131
rect 10652 4100 10977 4128
rect 10652 4088 10658 4100
rect 10965 4097 10977 4100
rect 11011 4097 11023 4131
rect 10965 4091 11023 4097
rect 14921 4131 14979 4137
rect 14921 4097 14933 4131
rect 14967 4128 14979 4131
rect 15286 4128 15292 4140
rect 14967 4100 15292 4128
rect 14967 4097 14979 4100
rect 14921 4091 14979 4097
rect 15286 4088 15292 4100
rect 15344 4088 15350 4140
rect 15654 4088 15660 4140
rect 15712 4088 15718 4140
rect 10686 4060 10692 4072
rect 10520 4032 10692 4060
rect 10229 4023 10287 4029
rect 10244 3992 10272 4023
rect 10686 4020 10692 4032
rect 10744 4020 10750 4072
rect 11057 4063 11115 4069
rect 11057 4029 11069 4063
rect 11103 4029 11115 4063
rect 11057 4023 11115 4029
rect 11072 3992 11100 4023
rect 11882 4020 11888 4072
rect 11940 4060 11946 4072
rect 12069 4063 12127 4069
rect 12069 4060 12081 4063
rect 11940 4032 12081 4060
rect 11940 4020 11946 4032
rect 12069 4029 12081 4032
rect 12115 4029 12127 4063
rect 12069 4023 12127 4029
rect 14737 4063 14795 4069
rect 14737 4029 14749 4063
rect 14783 4029 14795 4063
rect 15672 4060 15700 4088
rect 15933 4063 15991 4069
rect 15933 4060 15945 4063
rect 15672 4032 15945 4060
rect 14737 4023 14795 4029
rect 15933 4029 15945 4032
rect 15979 4029 15991 4063
rect 15933 4023 15991 4029
rect 16025 4063 16083 4069
rect 16025 4029 16037 4063
rect 16071 4029 16083 4063
rect 16025 4023 16083 4029
rect 14642 3992 14648 4004
rect 10244 3964 14648 3992
rect 14642 3952 14648 3964
rect 14700 3992 14706 4004
rect 14752 3992 14780 4023
rect 16040 3992 16068 4023
rect 14700 3964 16068 3992
rect 14700 3952 14706 3964
rect 9674 3884 9680 3936
rect 9732 3884 9738 3936
rect 10042 3884 10048 3936
rect 10100 3924 10106 3936
rect 10505 3927 10563 3933
rect 10505 3924 10517 3927
rect 10100 3896 10517 3924
rect 10100 3884 10106 3896
rect 10505 3893 10517 3896
rect 10551 3893 10563 3927
rect 10505 3887 10563 3893
rect 15378 3884 15384 3936
rect 15436 3884 15442 3936
rect 15473 3927 15531 3933
rect 15473 3893 15485 3927
rect 15519 3924 15531 3927
rect 15562 3924 15568 3936
rect 15519 3896 15568 3924
rect 15519 3893 15531 3896
rect 15473 3887 15531 3893
rect 15562 3884 15568 3896
rect 15620 3884 15626 3936
rect 1104 3834 31832 3856
rect 1104 3782 4182 3834
rect 4234 3782 4246 3834
rect 4298 3782 4310 3834
rect 4362 3782 4374 3834
rect 4426 3782 4438 3834
rect 4490 3782 4502 3834
rect 4554 3782 10182 3834
rect 10234 3782 10246 3834
rect 10298 3782 10310 3834
rect 10362 3782 10374 3834
rect 10426 3782 10438 3834
rect 10490 3782 10502 3834
rect 10554 3782 16182 3834
rect 16234 3782 16246 3834
rect 16298 3782 16310 3834
rect 16362 3782 16374 3834
rect 16426 3782 16438 3834
rect 16490 3782 16502 3834
rect 16554 3782 22182 3834
rect 22234 3782 22246 3834
rect 22298 3782 22310 3834
rect 22362 3782 22374 3834
rect 22426 3782 22438 3834
rect 22490 3782 22502 3834
rect 22554 3782 28182 3834
rect 28234 3782 28246 3834
rect 28298 3782 28310 3834
rect 28362 3782 28374 3834
rect 28426 3782 28438 3834
rect 28490 3782 28502 3834
rect 28554 3782 31832 3834
rect 1104 3760 31832 3782
rect 9674 3680 9680 3732
rect 9732 3680 9738 3732
rect 10042 3680 10048 3732
rect 10100 3680 10106 3732
rect 15378 3720 15384 3732
rect 15120 3692 15384 3720
rect 9692 3525 9720 3680
rect 9677 3519 9735 3525
rect 9677 3485 9689 3519
rect 9723 3485 9735 3519
rect 9677 3479 9735 3485
rect 9766 3476 9772 3528
rect 9824 3516 9830 3528
rect 10060 3525 10088 3680
rect 12158 3544 12164 3596
rect 12216 3544 12222 3596
rect 14550 3544 14556 3596
rect 14608 3544 14614 3596
rect 14642 3544 14648 3596
rect 14700 3544 14706 3596
rect 15120 3525 15148 3692
rect 15378 3680 15384 3692
rect 15436 3680 15442 3732
rect 15562 3680 15568 3732
rect 15620 3680 15626 3732
rect 17402 3680 17408 3732
rect 17460 3720 17466 3732
rect 17862 3720 17868 3732
rect 17460 3692 17868 3720
rect 17460 3680 17466 3692
rect 17862 3680 17868 3692
rect 17920 3680 17926 3732
rect 15194 3612 15200 3664
rect 15252 3652 15258 3664
rect 15289 3655 15347 3661
rect 15289 3652 15301 3655
rect 15252 3624 15301 3652
rect 15252 3612 15258 3624
rect 15289 3621 15301 3624
rect 15335 3621 15347 3655
rect 15580 3652 15608 3680
rect 15289 3615 15347 3621
rect 15396 3624 15608 3652
rect 15396 3525 15424 3624
rect 15470 3544 15476 3596
rect 15528 3584 15534 3596
rect 15657 3587 15715 3593
rect 15657 3584 15669 3587
rect 15528 3556 15669 3584
rect 15528 3544 15534 3556
rect 15657 3553 15669 3556
rect 15703 3553 15715 3587
rect 15657 3547 15715 3553
rect 9953 3519 10011 3525
rect 9953 3516 9965 3519
rect 9824 3488 9965 3516
rect 9824 3476 9830 3488
rect 9953 3485 9965 3488
rect 9999 3485 10011 3519
rect 9953 3479 10011 3485
rect 10045 3519 10103 3525
rect 10045 3485 10057 3519
rect 10091 3485 10103 3519
rect 10045 3479 10103 3485
rect 10321 3519 10379 3525
rect 10321 3485 10333 3519
rect 10367 3485 10379 3519
rect 10321 3479 10379 3485
rect 15105 3519 15163 3525
rect 15105 3485 15117 3519
rect 15151 3485 15163 3519
rect 15105 3479 15163 3485
rect 15381 3519 15439 3525
rect 15381 3485 15393 3519
rect 15427 3485 15439 3519
rect 15381 3479 15439 3485
rect 9030 3408 9036 3460
rect 9088 3448 9094 3460
rect 10336 3448 10364 3479
rect 9088 3420 10364 3448
rect 10597 3451 10655 3457
rect 9088 3408 9094 3420
rect 10597 3417 10609 3451
rect 10643 3417 10655 3451
rect 10597 3411 10655 3417
rect 9490 3340 9496 3392
rect 9548 3340 9554 3392
rect 9858 3340 9864 3392
rect 9916 3340 9922 3392
rect 10229 3383 10287 3389
rect 10229 3349 10241 3383
rect 10275 3380 10287 3383
rect 10612 3380 10640 3411
rect 11606 3408 11612 3460
rect 11664 3408 11670 3460
rect 12434 3408 12440 3460
rect 12492 3408 12498 3460
rect 13722 3448 13728 3460
rect 13662 3420 13728 3448
rect 13722 3408 13728 3420
rect 13780 3408 13786 3460
rect 14461 3451 14519 3457
rect 14461 3448 14473 3451
rect 13924 3420 14473 3448
rect 13924 3392 13952 3420
rect 14461 3417 14473 3420
rect 14507 3417 14519 3451
rect 14461 3411 14519 3417
rect 15933 3451 15991 3457
rect 15933 3417 15945 3451
rect 15979 3417 15991 3451
rect 15933 3411 15991 3417
rect 10275 3352 10640 3380
rect 10275 3349 10287 3352
rect 10229 3343 10287 3349
rect 11882 3340 11888 3392
rect 11940 3380 11946 3392
rect 12069 3383 12127 3389
rect 12069 3380 12081 3383
rect 11940 3352 12081 3380
rect 11940 3340 11946 3352
rect 12069 3349 12081 3352
rect 12115 3349 12127 3383
rect 12069 3343 12127 3349
rect 13906 3340 13912 3392
rect 13964 3340 13970 3392
rect 14090 3340 14096 3392
rect 14148 3340 14154 3392
rect 15565 3383 15623 3389
rect 15565 3349 15577 3383
rect 15611 3380 15623 3383
rect 15948 3380 15976 3411
rect 16666 3408 16672 3460
rect 16724 3408 16730 3460
rect 15611 3352 15976 3380
rect 15611 3349 15623 3352
rect 15565 3343 15623 3349
rect 1104 3290 31832 3312
rect 1104 3238 4922 3290
rect 4974 3238 4986 3290
rect 5038 3238 5050 3290
rect 5102 3238 5114 3290
rect 5166 3238 5178 3290
rect 5230 3238 5242 3290
rect 5294 3238 10922 3290
rect 10974 3238 10986 3290
rect 11038 3238 11050 3290
rect 11102 3238 11114 3290
rect 11166 3238 11178 3290
rect 11230 3238 11242 3290
rect 11294 3238 16922 3290
rect 16974 3238 16986 3290
rect 17038 3238 17050 3290
rect 17102 3238 17114 3290
rect 17166 3238 17178 3290
rect 17230 3238 17242 3290
rect 17294 3238 22922 3290
rect 22974 3238 22986 3290
rect 23038 3238 23050 3290
rect 23102 3238 23114 3290
rect 23166 3238 23178 3290
rect 23230 3238 23242 3290
rect 23294 3238 28922 3290
rect 28974 3238 28986 3290
rect 29038 3238 29050 3290
rect 29102 3238 29114 3290
rect 29166 3238 29178 3290
rect 29230 3238 29242 3290
rect 29294 3238 31832 3290
rect 1104 3216 31832 3238
rect 9490 3136 9496 3188
rect 9548 3136 9554 3188
rect 10778 3136 10784 3188
rect 10836 3136 10842 3188
rect 11606 3136 11612 3188
rect 11664 3136 11670 3188
rect 12434 3136 12440 3188
rect 12492 3176 12498 3188
rect 13081 3179 13139 3185
rect 13081 3176 13093 3179
rect 12492 3148 13093 3176
rect 12492 3136 12498 3148
rect 13081 3145 13093 3148
rect 13127 3145 13139 3179
rect 13081 3139 13139 3145
rect 13722 3136 13728 3188
rect 13780 3136 13786 3188
rect 14090 3136 14096 3188
rect 14148 3136 14154 3188
rect 16301 3179 16359 3185
rect 16301 3145 16313 3179
rect 16347 3176 16359 3179
rect 16574 3176 16580 3188
rect 16347 3148 16580 3176
rect 16347 3145 16359 3148
rect 16301 3139 16359 3145
rect 16574 3136 16580 3148
rect 16632 3136 16638 3188
rect 16666 3136 16672 3188
rect 16724 3176 16730 3188
rect 16761 3179 16819 3185
rect 16761 3176 16773 3179
rect 16724 3148 16773 3176
rect 16724 3136 16730 3148
rect 16761 3145 16773 3148
rect 16807 3145 16819 3179
rect 16761 3139 16819 3145
rect 9309 3111 9367 3117
rect 9309 3077 9321 3111
rect 9355 3108 9367 3111
rect 9508 3108 9536 3136
rect 9355 3080 9536 3108
rect 9355 3077 9367 3080
rect 9309 3071 9367 3077
rect 9858 3068 9864 3120
rect 9916 3068 9922 3120
rect 14108 3108 14136 3136
rect 13280 3080 14136 3108
rect 6914 3000 6920 3052
rect 6972 3040 6978 3052
rect 9030 3040 9036 3052
rect 6972 3012 9036 3040
rect 6972 3000 6978 3012
rect 9030 3000 9036 3012
rect 9088 3000 9094 3052
rect 13280 3049 13308 3080
rect 11701 3043 11759 3049
rect 11701 3009 11713 3043
rect 11747 3009 11759 3043
rect 11701 3003 11759 3009
rect 13265 3043 13323 3049
rect 13265 3009 13277 3043
rect 13311 3009 13323 3043
rect 13265 3003 13323 3009
rect 13817 3043 13875 3049
rect 13817 3009 13829 3043
rect 13863 3040 13875 3043
rect 16209 3043 16267 3049
rect 16209 3040 16221 3043
rect 13863 3012 16221 3040
rect 13863 3009 13875 3012
rect 13817 3003 13875 3009
rect 16209 3009 16221 3012
rect 16255 3040 16267 3043
rect 16669 3043 16727 3049
rect 16669 3040 16681 3043
rect 16255 3012 16681 3040
rect 16255 3009 16267 3012
rect 16209 3003 16267 3009
rect 16669 3009 16681 3012
rect 16715 3009 16727 3043
rect 16669 3003 16727 3009
rect 9766 2932 9772 2984
rect 9824 2972 9830 2984
rect 11716 2972 11744 3003
rect 13832 2972 13860 3003
rect 9824 2944 13860 2972
rect 9824 2932 9830 2944
rect 1104 2746 31832 2768
rect 1104 2694 4182 2746
rect 4234 2694 4246 2746
rect 4298 2694 4310 2746
rect 4362 2694 4374 2746
rect 4426 2694 4438 2746
rect 4490 2694 4502 2746
rect 4554 2694 10182 2746
rect 10234 2694 10246 2746
rect 10298 2694 10310 2746
rect 10362 2694 10374 2746
rect 10426 2694 10438 2746
rect 10490 2694 10502 2746
rect 10554 2694 16182 2746
rect 16234 2694 16246 2746
rect 16298 2694 16310 2746
rect 16362 2694 16374 2746
rect 16426 2694 16438 2746
rect 16490 2694 16502 2746
rect 16554 2694 22182 2746
rect 22234 2694 22246 2746
rect 22298 2694 22310 2746
rect 22362 2694 22374 2746
rect 22426 2694 22438 2746
rect 22490 2694 22502 2746
rect 22554 2694 28182 2746
rect 28234 2694 28246 2746
rect 28298 2694 28310 2746
rect 28362 2694 28374 2746
rect 28426 2694 28438 2746
rect 28490 2694 28502 2746
rect 28554 2694 31832 2746
rect 1104 2672 31832 2694
rect 29273 2635 29331 2641
rect 29273 2601 29285 2635
rect 29319 2632 29331 2635
rect 29362 2632 29368 2644
rect 29319 2604 29368 2632
rect 29319 2601 29331 2604
rect 29273 2595 29331 2601
rect 29362 2592 29368 2604
rect 29420 2592 29426 2644
rect 13906 2496 13912 2508
rect 6886 2468 13912 2496
rect 1765 2431 1823 2437
rect 1765 2397 1777 2431
rect 1811 2428 1823 2431
rect 6886 2428 6914 2468
rect 13906 2456 13912 2468
rect 13964 2456 13970 2508
rect 1811 2400 6914 2428
rect 1811 2397 1823 2400
rect 1765 2391 1823 2397
rect 11882 2388 11888 2440
rect 11940 2388 11946 2440
rect 17034 2388 17040 2440
rect 17092 2428 17098 2440
rect 17589 2431 17647 2437
rect 17589 2428 17601 2431
rect 17092 2400 17601 2428
rect 17092 2388 17098 2400
rect 17589 2397 17601 2400
rect 17635 2397 17647 2431
rect 17589 2391 17647 2397
rect 17862 2388 17868 2440
rect 17920 2428 17926 2440
rect 23385 2431 23443 2437
rect 23385 2428 23397 2431
rect 17920 2400 23397 2428
rect 17920 2388 17926 2400
rect 23385 2397 23397 2400
rect 23431 2397 23443 2431
rect 23385 2391 23443 2397
rect 29089 2431 29147 2437
rect 29089 2397 29101 2431
rect 29135 2428 29147 2431
rect 29362 2428 29368 2440
rect 29135 2400 29368 2428
rect 29135 2397 29147 2400
rect 29089 2391 29147 2397
rect 29362 2388 29368 2400
rect 29420 2388 29426 2440
rect 31202 2388 31208 2440
rect 31260 2388 31266 2440
rect 14 2320 20 2372
rect 72 2360 78 2372
rect 1397 2363 1455 2369
rect 1397 2360 1409 2363
rect 72 2332 1409 2360
rect 72 2320 78 2332
rect 1397 2329 1409 2332
rect 1443 2329 1455 2363
rect 1397 2323 1455 2329
rect 6089 2363 6147 2369
rect 6089 2329 6101 2363
rect 6135 2360 6147 2363
rect 10778 2360 10784 2372
rect 6135 2332 10784 2360
rect 6135 2329 6147 2332
rect 6089 2323 6147 2329
rect 10778 2320 10784 2332
rect 10836 2320 10842 2372
rect 5810 2252 5816 2304
rect 5868 2252 5874 2304
rect 11606 2252 11612 2304
rect 11664 2252 11670 2304
rect 17402 2252 17408 2304
rect 17460 2292 17466 2304
rect 17681 2295 17739 2301
rect 17681 2292 17693 2295
rect 17460 2264 17693 2292
rect 17460 2252 17466 2264
rect 17681 2261 17693 2264
rect 17727 2261 17739 2295
rect 17681 2255 17739 2261
rect 23474 2252 23480 2304
rect 23532 2252 23538 2304
rect 31386 2252 31392 2304
rect 31444 2252 31450 2304
rect 1104 2202 31832 2224
rect 1104 2150 4922 2202
rect 4974 2150 4986 2202
rect 5038 2150 5050 2202
rect 5102 2150 5114 2202
rect 5166 2150 5178 2202
rect 5230 2150 5242 2202
rect 5294 2150 10922 2202
rect 10974 2150 10986 2202
rect 11038 2150 11050 2202
rect 11102 2150 11114 2202
rect 11166 2150 11178 2202
rect 11230 2150 11242 2202
rect 11294 2150 16922 2202
rect 16974 2150 16986 2202
rect 17038 2150 17050 2202
rect 17102 2150 17114 2202
rect 17166 2150 17178 2202
rect 17230 2150 17242 2202
rect 17294 2150 22922 2202
rect 22974 2150 22986 2202
rect 23038 2150 23050 2202
rect 23102 2150 23114 2202
rect 23166 2150 23178 2202
rect 23230 2150 23242 2202
rect 23294 2150 28922 2202
rect 28974 2150 28986 2202
rect 29038 2150 29050 2202
rect 29102 2150 29114 2202
rect 29166 2150 29178 2202
rect 29230 2150 29242 2202
rect 29294 2150 31832 2202
rect 1104 2128 31832 2150
<< via1 >>
rect 4922 32614 4974 32666
rect 4986 32614 5038 32666
rect 5050 32614 5102 32666
rect 5114 32614 5166 32666
rect 5178 32614 5230 32666
rect 5242 32614 5294 32666
rect 10922 32614 10974 32666
rect 10986 32614 11038 32666
rect 11050 32614 11102 32666
rect 11114 32614 11166 32666
rect 11178 32614 11230 32666
rect 11242 32614 11294 32666
rect 16922 32614 16974 32666
rect 16986 32614 17038 32666
rect 17050 32614 17102 32666
rect 17114 32614 17166 32666
rect 17178 32614 17230 32666
rect 17242 32614 17294 32666
rect 22922 32614 22974 32666
rect 22986 32614 23038 32666
rect 23050 32614 23102 32666
rect 23114 32614 23166 32666
rect 23178 32614 23230 32666
rect 23242 32614 23294 32666
rect 28922 32614 28974 32666
rect 28986 32614 29038 32666
rect 29050 32614 29102 32666
rect 29114 32614 29166 32666
rect 29178 32614 29230 32666
rect 29242 32614 29294 32666
rect 1308 32512 1360 32564
rect 18696 32512 18748 32564
rect 24492 32512 24544 32564
rect 7104 32376 7156 32428
rect 12900 32376 12952 32428
rect 19340 32419 19392 32428
rect 19340 32385 19349 32419
rect 19349 32385 19383 32419
rect 19383 32385 19392 32419
rect 19340 32376 19392 32385
rect 24676 32419 24728 32428
rect 24676 32385 24685 32419
rect 24685 32385 24719 32419
rect 24719 32385 24728 32419
rect 24676 32376 24728 32385
rect 30288 32376 30340 32428
rect 12440 32240 12492 32292
rect 7380 32215 7432 32224
rect 7380 32181 7389 32215
rect 7389 32181 7423 32215
rect 7423 32181 7432 32215
rect 7380 32172 7432 32181
rect 13176 32215 13228 32224
rect 13176 32181 13185 32215
rect 13185 32181 13219 32215
rect 13219 32181 13228 32215
rect 13176 32172 13228 32181
rect 30564 32215 30616 32224
rect 30564 32181 30573 32215
rect 30573 32181 30607 32215
rect 30607 32181 30616 32215
rect 30564 32172 30616 32181
rect 4182 32070 4234 32122
rect 4246 32070 4298 32122
rect 4310 32070 4362 32122
rect 4374 32070 4426 32122
rect 4438 32070 4490 32122
rect 4502 32070 4554 32122
rect 10182 32070 10234 32122
rect 10246 32070 10298 32122
rect 10310 32070 10362 32122
rect 10374 32070 10426 32122
rect 10438 32070 10490 32122
rect 10502 32070 10554 32122
rect 16182 32070 16234 32122
rect 16246 32070 16298 32122
rect 16310 32070 16362 32122
rect 16374 32070 16426 32122
rect 16438 32070 16490 32122
rect 16502 32070 16554 32122
rect 22182 32070 22234 32122
rect 22246 32070 22298 32122
rect 22310 32070 22362 32122
rect 22374 32070 22426 32122
rect 22438 32070 22490 32122
rect 22502 32070 22554 32122
rect 28182 32070 28234 32122
rect 28246 32070 28298 32122
rect 28310 32070 28362 32122
rect 28374 32070 28426 32122
rect 28438 32070 28490 32122
rect 28502 32070 28554 32122
rect 20168 31764 20220 31816
rect 13544 31696 13596 31748
rect 18236 31628 18288 31680
rect 19340 31628 19392 31680
rect 4922 31526 4974 31578
rect 4986 31526 5038 31578
rect 5050 31526 5102 31578
rect 5114 31526 5166 31578
rect 5178 31526 5230 31578
rect 5242 31526 5294 31578
rect 10922 31526 10974 31578
rect 10986 31526 11038 31578
rect 11050 31526 11102 31578
rect 11114 31526 11166 31578
rect 11178 31526 11230 31578
rect 11242 31526 11294 31578
rect 16922 31526 16974 31578
rect 16986 31526 17038 31578
rect 17050 31526 17102 31578
rect 17114 31526 17166 31578
rect 17178 31526 17230 31578
rect 17242 31526 17294 31578
rect 22922 31526 22974 31578
rect 22986 31526 23038 31578
rect 23050 31526 23102 31578
rect 23114 31526 23166 31578
rect 23178 31526 23230 31578
rect 23242 31526 23294 31578
rect 28922 31526 28974 31578
rect 28986 31526 29038 31578
rect 29050 31526 29102 31578
rect 29114 31526 29166 31578
rect 29178 31526 29230 31578
rect 29242 31526 29294 31578
rect 13544 31467 13596 31476
rect 13544 31433 13553 31467
rect 13553 31433 13587 31467
rect 13587 31433 13596 31467
rect 13544 31424 13596 31433
rect 24676 31424 24728 31476
rect 14004 31356 14056 31408
rect 14372 31356 14424 31408
rect 14832 31356 14884 31408
rect 16764 31288 16816 31340
rect 10784 31220 10836 31272
rect 12808 31220 12860 31272
rect 12900 31263 12952 31272
rect 12900 31229 12909 31263
rect 12909 31229 12943 31263
rect 12943 31229 12952 31263
rect 12900 31220 12952 31229
rect 14096 31263 14148 31272
rect 14096 31229 14105 31263
rect 14105 31229 14139 31263
rect 14139 31229 14148 31263
rect 14096 31220 14148 31229
rect 17224 31288 17276 31340
rect 17500 31331 17552 31340
rect 17500 31297 17509 31331
rect 17509 31297 17543 31331
rect 17543 31297 17552 31331
rect 17500 31288 17552 31297
rect 18236 31356 18288 31408
rect 17868 31331 17920 31340
rect 17868 31297 17877 31331
rect 17877 31297 17911 31331
rect 17911 31297 17920 31331
rect 17868 31288 17920 31297
rect 17592 31220 17644 31272
rect 19432 31356 19484 31408
rect 18788 31220 18840 31272
rect 11612 31127 11664 31136
rect 11612 31093 11621 31127
rect 11621 31093 11655 31127
rect 11655 31093 11664 31127
rect 11612 31084 11664 31093
rect 13176 31127 13228 31136
rect 13176 31093 13185 31127
rect 13185 31093 13219 31127
rect 13219 31093 13228 31127
rect 13176 31084 13228 31093
rect 15476 31084 15528 31136
rect 16856 31127 16908 31136
rect 16856 31093 16865 31127
rect 16865 31093 16899 31127
rect 16899 31093 16908 31127
rect 16856 31084 16908 31093
rect 17316 31127 17368 31136
rect 17316 31093 17325 31127
rect 17325 31093 17359 31127
rect 17359 31093 17368 31127
rect 17316 31084 17368 31093
rect 20168 31195 20220 31204
rect 20168 31161 20177 31195
rect 20177 31161 20211 31195
rect 20211 31161 20220 31195
rect 20168 31152 20220 31161
rect 17776 31084 17828 31136
rect 18512 31084 18564 31136
rect 4182 30982 4234 31034
rect 4246 30982 4298 31034
rect 4310 30982 4362 31034
rect 4374 30982 4426 31034
rect 4438 30982 4490 31034
rect 4502 30982 4554 31034
rect 10182 30982 10234 31034
rect 10246 30982 10298 31034
rect 10310 30982 10362 31034
rect 10374 30982 10426 31034
rect 10438 30982 10490 31034
rect 10502 30982 10554 31034
rect 16182 30982 16234 31034
rect 16246 30982 16298 31034
rect 16310 30982 16362 31034
rect 16374 30982 16426 31034
rect 16438 30982 16490 31034
rect 16502 30982 16554 31034
rect 22182 30982 22234 31034
rect 22246 30982 22298 31034
rect 22310 30982 22362 31034
rect 22374 30982 22426 31034
rect 22438 30982 22490 31034
rect 22502 30982 22554 31034
rect 28182 30982 28234 31034
rect 28246 30982 28298 31034
rect 28310 30982 28362 31034
rect 28374 30982 28426 31034
rect 28438 30982 28490 31034
rect 28502 30982 28554 31034
rect 11612 30744 11664 30796
rect 13176 30880 13228 30932
rect 13544 30880 13596 30932
rect 14096 30880 14148 30932
rect 14832 30923 14884 30932
rect 14832 30889 14841 30923
rect 14841 30889 14875 30923
rect 14875 30889 14884 30923
rect 14832 30880 14884 30889
rect 17316 30880 17368 30932
rect 17592 30880 17644 30932
rect 12900 30812 12952 30864
rect 940 30676 992 30728
rect 10784 30719 10836 30728
rect 10784 30685 10793 30719
rect 10793 30685 10827 30719
rect 10827 30685 10836 30719
rect 10784 30676 10836 30685
rect 12440 30676 12492 30728
rect 12992 30676 13044 30728
rect 15476 30787 15528 30796
rect 15476 30753 15485 30787
rect 15485 30753 15519 30787
rect 15519 30753 15528 30787
rect 15476 30744 15528 30753
rect 1584 30583 1636 30592
rect 1584 30549 1593 30583
rect 1593 30549 1627 30583
rect 1627 30549 1636 30583
rect 1584 30540 1636 30549
rect 13452 30651 13504 30660
rect 13452 30617 13461 30651
rect 13461 30617 13495 30651
rect 13495 30617 13504 30651
rect 13452 30608 13504 30617
rect 14096 30608 14148 30660
rect 15016 30676 15068 30728
rect 16856 30676 16908 30728
rect 15752 30651 15804 30660
rect 15752 30617 15761 30651
rect 15761 30617 15795 30651
rect 15795 30617 15804 30651
rect 15752 30608 15804 30617
rect 14188 30583 14240 30592
rect 14188 30549 14197 30583
rect 14197 30549 14231 30583
rect 14231 30549 14240 30583
rect 14188 30540 14240 30549
rect 14280 30540 14332 30592
rect 14372 30540 14424 30592
rect 16580 30540 16632 30592
rect 18144 30719 18196 30728
rect 18144 30685 18153 30719
rect 18153 30685 18187 30719
rect 18187 30685 18196 30719
rect 18144 30676 18196 30685
rect 18788 30676 18840 30728
rect 17316 30608 17368 30660
rect 17868 30608 17920 30660
rect 17408 30583 17460 30592
rect 17408 30549 17417 30583
rect 17417 30549 17451 30583
rect 17451 30549 17460 30583
rect 17408 30540 17460 30549
rect 17592 30540 17644 30592
rect 19340 30676 19392 30728
rect 19524 30608 19576 30660
rect 4922 30438 4974 30490
rect 4986 30438 5038 30490
rect 5050 30438 5102 30490
rect 5114 30438 5166 30490
rect 5178 30438 5230 30490
rect 5242 30438 5294 30490
rect 10922 30438 10974 30490
rect 10986 30438 11038 30490
rect 11050 30438 11102 30490
rect 11114 30438 11166 30490
rect 11178 30438 11230 30490
rect 11242 30438 11294 30490
rect 16922 30438 16974 30490
rect 16986 30438 17038 30490
rect 17050 30438 17102 30490
rect 17114 30438 17166 30490
rect 17178 30438 17230 30490
rect 17242 30438 17294 30490
rect 22922 30438 22974 30490
rect 22986 30438 23038 30490
rect 23050 30438 23102 30490
rect 23114 30438 23166 30490
rect 23178 30438 23230 30490
rect 23242 30438 23294 30490
rect 28922 30438 28974 30490
rect 28986 30438 29038 30490
rect 29050 30438 29102 30490
rect 29114 30438 29166 30490
rect 29178 30438 29230 30490
rect 29242 30438 29294 30490
rect 12808 30336 12860 30388
rect 15752 30336 15804 30388
rect 11888 30243 11940 30252
rect 11888 30209 11897 30243
rect 11897 30209 11931 30243
rect 11931 30209 11940 30243
rect 11888 30200 11940 30209
rect 12900 30200 12952 30252
rect 13912 30243 13964 30252
rect 13912 30209 13921 30243
rect 13921 30209 13955 30243
rect 13955 30209 13964 30243
rect 13912 30200 13964 30209
rect 14924 30243 14976 30252
rect 14924 30209 14933 30243
rect 14933 30209 14967 30243
rect 14967 30209 14976 30243
rect 14924 30200 14976 30209
rect 15016 30200 15068 30252
rect 14648 30132 14700 30184
rect 13636 29996 13688 30048
rect 14096 29996 14148 30048
rect 15752 30243 15804 30252
rect 15752 30209 15794 30243
rect 15794 30209 15804 30243
rect 15752 30200 15804 30209
rect 16672 30268 16724 30320
rect 17408 30200 17460 30252
rect 17500 30200 17552 30252
rect 17776 30200 17828 30252
rect 18144 30200 18196 30252
rect 19708 30268 19760 30320
rect 18512 30243 18564 30252
rect 18512 30209 18521 30243
rect 18521 30209 18555 30243
rect 18555 30209 18564 30243
rect 18512 30200 18564 30209
rect 18788 30175 18840 30184
rect 16764 29996 16816 30048
rect 16856 29996 16908 30048
rect 17960 29996 18012 30048
rect 18788 30141 18797 30175
rect 18797 30141 18831 30175
rect 18831 30141 18840 30175
rect 18788 30132 18840 30141
rect 19524 30132 19576 30184
rect 20444 29996 20496 30048
rect 4182 29894 4234 29946
rect 4246 29894 4298 29946
rect 4310 29894 4362 29946
rect 4374 29894 4426 29946
rect 4438 29894 4490 29946
rect 4502 29894 4554 29946
rect 10182 29894 10234 29946
rect 10246 29894 10298 29946
rect 10310 29894 10362 29946
rect 10374 29894 10426 29946
rect 10438 29894 10490 29946
rect 10502 29894 10554 29946
rect 16182 29894 16234 29946
rect 16246 29894 16298 29946
rect 16310 29894 16362 29946
rect 16374 29894 16426 29946
rect 16438 29894 16490 29946
rect 16502 29894 16554 29946
rect 22182 29894 22234 29946
rect 22246 29894 22298 29946
rect 22310 29894 22362 29946
rect 22374 29894 22426 29946
rect 22438 29894 22490 29946
rect 22502 29894 22554 29946
rect 28182 29894 28234 29946
rect 28246 29894 28298 29946
rect 28310 29894 28362 29946
rect 28374 29894 28426 29946
rect 28438 29894 28490 29946
rect 28502 29894 28554 29946
rect 13912 29835 13964 29844
rect 13912 29801 13921 29835
rect 13921 29801 13955 29835
rect 13955 29801 13964 29835
rect 13912 29792 13964 29801
rect 14004 29792 14056 29844
rect 14924 29792 14976 29844
rect 16672 29835 16724 29844
rect 16672 29801 16681 29835
rect 16681 29801 16715 29835
rect 16715 29801 16724 29835
rect 16672 29792 16724 29801
rect 16764 29792 16816 29844
rect 17408 29792 17460 29844
rect 17500 29792 17552 29844
rect 19432 29835 19484 29844
rect 19432 29801 19441 29835
rect 19441 29801 19475 29835
rect 19475 29801 19484 29835
rect 19432 29792 19484 29801
rect 19708 29835 19760 29844
rect 19708 29801 19717 29835
rect 19717 29801 19751 29835
rect 19751 29801 19760 29835
rect 19708 29792 19760 29801
rect 12992 29699 13044 29708
rect 12992 29665 13001 29699
rect 13001 29665 13035 29699
rect 13035 29665 13044 29699
rect 12992 29656 13044 29665
rect 14188 29588 14240 29640
rect 14280 29631 14332 29640
rect 14280 29597 14289 29631
rect 14289 29597 14323 29631
rect 14323 29597 14332 29631
rect 14280 29588 14332 29597
rect 16028 29724 16080 29776
rect 16580 29631 16632 29640
rect 16580 29597 16589 29631
rect 16589 29597 16623 29631
rect 16623 29597 16632 29631
rect 16580 29588 16632 29597
rect 17500 29699 17552 29708
rect 17500 29665 17509 29699
rect 17509 29665 17543 29699
rect 17543 29665 17552 29699
rect 17500 29656 17552 29665
rect 18512 29656 18564 29708
rect 17592 29520 17644 29572
rect 18052 29588 18104 29640
rect 20444 29588 20496 29640
rect 13268 29495 13320 29504
rect 13268 29461 13277 29495
rect 13277 29461 13311 29495
rect 13311 29461 13320 29495
rect 13268 29452 13320 29461
rect 13636 29452 13688 29504
rect 15016 29452 15068 29504
rect 15752 29452 15804 29504
rect 16856 29495 16908 29504
rect 16856 29461 16873 29495
rect 16873 29461 16908 29495
rect 16856 29452 16908 29461
rect 17408 29452 17460 29504
rect 4922 29350 4974 29402
rect 4986 29350 5038 29402
rect 5050 29350 5102 29402
rect 5114 29350 5166 29402
rect 5178 29350 5230 29402
rect 5242 29350 5294 29402
rect 10922 29350 10974 29402
rect 10986 29350 11038 29402
rect 11050 29350 11102 29402
rect 11114 29350 11166 29402
rect 11178 29350 11230 29402
rect 11242 29350 11294 29402
rect 16922 29350 16974 29402
rect 16986 29350 17038 29402
rect 17050 29350 17102 29402
rect 17114 29350 17166 29402
rect 17178 29350 17230 29402
rect 17242 29350 17294 29402
rect 22922 29350 22974 29402
rect 22986 29350 23038 29402
rect 23050 29350 23102 29402
rect 23114 29350 23166 29402
rect 23178 29350 23230 29402
rect 23242 29350 23294 29402
rect 28922 29350 28974 29402
rect 28986 29350 29038 29402
rect 29050 29350 29102 29402
rect 29114 29350 29166 29402
rect 29178 29350 29230 29402
rect 29242 29350 29294 29402
rect 13268 29112 13320 29164
rect 13728 29112 13780 29164
rect 14372 29112 14424 29164
rect 15752 29044 15804 29096
rect 4182 28806 4234 28858
rect 4246 28806 4298 28858
rect 4310 28806 4362 28858
rect 4374 28806 4426 28858
rect 4438 28806 4490 28858
rect 4502 28806 4554 28858
rect 10182 28806 10234 28858
rect 10246 28806 10298 28858
rect 10310 28806 10362 28858
rect 10374 28806 10426 28858
rect 10438 28806 10490 28858
rect 10502 28806 10554 28858
rect 16182 28806 16234 28858
rect 16246 28806 16298 28858
rect 16310 28806 16362 28858
rect 16374 28806 16426 28858
rect 16438 28806 16490 28858
rect 16502 28806 16554 28858
rect 22182 28806 22234 28858
rect 22246 28806 22298 28858
rect 22310 28806 22362 28858
rect 22374 28806 22426 28858
rect 22438 28806 22490 28858
rect 22502 28806 22554 28858
rect 28182 28806 28234 28858
rect 28246 28806 28298 28858
rect 28310 28806 28362 28858
rect 28374 28806 28426 28858
rect 28438 28806 28490 28858
rect 28502 28806 28554 28858
rect 11888 28704 11940 28756
rect 8484 28543 8536 28552
rect 8484 28509 8493 28543
rect 8493 28509 8527 28543
rect 8527 28509 8536 28543
rect 8484 28500 8536 28509
rect 8668 28500 8720 28552
rect 14372 28543 14424 28552
rect 14372 28509 14381 28543
rect 14381 28509 14415 28543
rect 14415 28509 14424 28543
rect 14372 28500 14424 28509
rect 10784 28432 10836 28484
rect 10324 28407 10376 28416
rect 10324 28373 10333 28407
rect 10333 28373 10367 28407
rect 10367 28373 10376 28407
rect 10324 28364 10376 28373
rect 10508 28364 10560 28416
rect 13820 28432 13872 28484
rect 14004 28364 14056 28416
rect 14096 28407 14148 28416
rect 14096 28373 14105 28407
rect 14105 28373 14139 28407
rect 14139 28373 14148 28407
rect 14096 28364 14148 28373
rect 14924 28500 14976 28552
rect 14740 28432 14792 28484
rect 14556 28364 14608 28416
rect 4922 28262 4974 28314
rect 4986 28262 5038 28314
rect 5050 28262 5102 28314
rect 5114 28262 5166 28314
rect 5178 28262 5230 28314
rect 5242 28262 5294 28314
rect 10922 28262 10974 28314
rect 10986 28262 11038 28314
rect 11050 28262 11102 28314
rect 11114 28262 11166 28314
rect 11178 28262 11230 28314
rect 11242 28262 11294 28314
rect 16922 28262 16974 28314
rect 16986 28262 17038 28314
rect 17050 28262 17102 28314
rect 17114 28262 17166 28314
rect 17178 28262 17230 28314
rect 17242 28262 17294 28314
rect 22922 28262 22974 28314
rect 22986 28262 23038 28314
rect 23050 28262 23102 28314
rect 23114 28262 23166 28314
rect 23178 28262 23230 28314
rect 23242 28262 23294 28314
rect 28922 28262 28974 28314
rect 28986 28262 29038 28314
rect 29050 28262 29102 28314
rect 29114 28262 29166 28314
rect 29178 28262 29230 28314
rect 29242 28262 29294 28314
rect 8484 28160 8536 28212
rect 10508 28160 10560 28212
rect 13728 28203 13780 28212
rect 13728 28169 13737 28203
rect 13737 28169 13771 28203
rect 13771 28169 13780 28203
rect 13728 28160 13780 28169
rect 13820 28203 13872 28212
rect 13820 28169 13829 28203
rect 13829 28169 13863 28203
rect 13863 28169 13872 28203
rect 13820 28160 13872 28169
rect 14096 28160 14148 28212
rect 14372 28160 14424 28212
rect 14464 28160 14516 28212
rect 9220 27999 9272 28008
rect 9220 27965 9229 27999
rect 9229 27965 9263 27999
rect 9263 27965 9272 27999
rect 9220 27956 9272 27965
rect 9864 27956 9916 28008
rect 10324 27999 10376 28008
rect 10324 27965 10333 27999
rect 10333 27965 10367 27999
rect 10367 27965 10376 27999
rect 10324 27956 10376 27965
rect 11888 28024 11940 28076
rect 13912 28024 13964 28076
rect 14280 28067 14332 28076
rect 14280 28033 14289 28067
rect 14289 28033 14323 28067
rect 14323 28033 14332 28067
rect 14280 28024 14332 28033
rect 14372 28067 14424 28076
rect 14372 28033 14381 28067
rect 14381 28033 14415 28067
rect 14415 28033 14424 28067
rect 14372 28024 14424 28033
rect 14648 28024 14700 28076
rect 10692 27956 10744 28008
rect 13728 27956 13780 28008
rect 7840 27820 7892 27872
rect 14004 27931 14056 27940
rect 14004 27897 14013 27931
rect 14013 27897 14047 27931
rect 14047 27897 14056 27931
rect 14004 27888 14056 27897
rect 14372 27888 14424 27940
rect 14740 27956 14792 28008
rect 17592 28092 17644 28144
rect 16580 27956 16632 28008
rect 18880 28024 18932 28076
rect 20352 28067 20404 28076
rect 20352 28033 20361 28067
rect 20361 28033 20395 28067
rect 20395 28033 20404 28067
rect 20352 28024 20404 28033
rect 23388 28067 23440 28076
rect 23388 28033 23397 28067
rect 23397 28033 23431 28067
rect 23431 28033 23440 28067
rect 23388 28024 23440 28033
rect 26608 28067 26660 28076
rect 26608 28033 26617 28067
rect 26617 28033 26651 28067
rect 26651 28033 26660 28067
rect 26608 28024 26660 28033
rect 11336 27820 11388 27872
rect 14096 27863 14148 27872
rect 14096 27829 14105 27863
rect 14105 27829 14139 27863
rect 14139 27829 14148 27863
rect 14096 27820 14148 27829
rect 14280 27820 14332 27872
rect 15844 27820 15896 27872
rect 16948 27956 17000 28008
rect 17684 27956 17736 28008
rect 18052 27999 18104 28008
rect 18052 27965 18061 27999
rect 18061 27965 18095 27999
rect 18095 27965 18104 27999
rect 18052 27956 18104 27965
rect 18972 27956 19024 28008
rect 20168 27956 20220 28008
rect 19984 27888 20036 27940
rect 20720 27931 20772 27940
rect 20720 27897 20729 27931
rect 20729 27897 20763 27931
rect 20763 27897 20772 27931
rect 20720 27888 20772 27897
rect 16672 27863 16724 27872
rect 16672 27829 16681 27863
rect 16681 27829 16715 27863
rect 16715 27829 16724 27863
rect 16672 27820 16724 27829
rect 16764 27820 16816 27872
rect 17776 27820 17828 27872
rect 23112 27820 23164 27872
rect 26332 27820 26384 27872
rect 4182 27718 4234 27770
rect 4246 27718 4298 27770
rect 4310 27718 4362 27770
rect 4374 27718 4426 27770
rect 4438 27718 4490 27770
rect 4502 27718 4554 27770
rect 10182 27718 10234 27770
rect 10246 27718 10298 27770
rect 10310 27718 10362 27770
rect 10374 27718 10426 27770
rect 10438 27718 10490 27770
rect 10502 27718 10554 27770
rect 16182 27718 16234 27770
rect 16246 27718 16298 27770
rect 16310 27718 16362 27770
rect 16374 27718 16426 27770
rect 16438 27718 16490 27770
rect 16502 27718 16554 27770
rect 22182 27718 22234 27770
rect 22246 27718 22298 27770
rect 22310 27718 22362 27770
rect 22374 27718 22426 27770
rect 22438 27718 22490 27770
rect 22502 27718 22554 27770
rect 28182 27718 28234 27770
rect 28246 27718 28298 27770
rect 28310 27718 28362 27770
rect 28374 27718 28426 27770
rect 28438 27718 28490 27770
rect 28502 27718 28554 27770
rect 14924 27616 14976 27668
rect 15568 27616 15620 27668
rect 16488 27616 16540 27668
rect 13912 27480 13964 27532
rect 8668 27412 8720 27464
rect 4804 27344 4856 27396
rect 9128 27344 9180 27396
rect 9312 27387 9364 27396
rect 9312 27353 9346 27387
rect 9346 27353 9364 27387
rect 9312 27344 9364 27353
rect 10048 27276 10100 27328
rect 14096 27412 14148 27464
rect 10600 27344 10652 27396
rect 14464 27480 14516 27532
rect 15016 27548 15068 27600
rect 16672 27548 16724 27600
rect 16948 27548 17000 27600
rect 17408 27591 17460 27600
rect 17408 27557 17417 27591
rect 17417 27557 17451 27591
rect 17451 27557 17460 27591
rect 17408 27548 17460 27557
rect 17868 27616 17920 27668
rect 18420 27616 18472 27668
rect 16028 27480 16080 27532
rect 18328 27548 18380 27600
rect 19708 27548 19760 27600
rect 29368 27548 29420 27600
rect 30564 27548 30616 27600
rect 15016 27412 15068 27464
rect 17868 27412 17920 27464
rect 18052 27455 18104 27464
rect 18052 27421 18061 27455
rect 18061 27421 18095 27455
rect 18095 27421 18104 27455
rect 18052 27412 18104 27421
rect 16764 27344 16816 27396
rect 17408 27344 17460 27396
rect 18328 27387 18380 27396
rect 18328 27353 18337 27387
rect 18337 27353 18371 27387
rect 18371 27353 18380 27387
rect 18328 27344 18380 27353
rect 18512 27412 18564 27464
rect 19340 27523 19392 27532
rect 19340 27489 19349 27523
rect 19349 27489 19383 27523
rect 19383 27489 19392 27523
rect 19340 27480 19392 27489
rect 19984 27523 20036 27532
rect 19984 27489 19993 27523
rect 19993 27489 20027 27523
rect 20027 27489 20036 27523
rect 19984 27480 20036 27489
rect 18972 27455 19024 27464
rect 18972 27421 18981 27455
rect 18981 27421 19015 27455
rect 19015 27421 19024 27455
rect 18972 27412 19024 27421
rect 19892 27412 19944 27464
rect 20076 27455 20128 27464
rect 20076 27421 20085 27455
rect 20085 27421 20119 27455
rect 20119 27421 20128 27455
rect 20076 27412 20128 27421
rect 20720 27412 20772 27464
rect 22836 27455 22888 27464
rect 22836 27421 22845 27455
rect 22845 27421 22879 27455
rect 22879 27421 22888 27455
rect 22836 27412 22888 27421
rect 23112 27455 23164 27464
rect 23112 27421 23146 27455
rect 23146 27421 23164 27455
rect 23112 27412 23164 27421
rect 25320 27412 25372 27464
rect 26332 27455 26384 27464
rect 26332 27421 26366 27455
rect 26366 27421 26384 27455
rect 26332 27412 26384 27421
rect 10508 27319 10560 27328
rect 10508 27285 10517 27319
rect 10517 27285 10551 27319
rect 10551 27285 10560 27319
rect 10508 27276 10560 27285
rect 14556 27319 14608 27328
rect 14556 27285 14565 27319
rect 14565 27285 14599 27319
rect 14599 27285 14608 27319
rect 14556 27276 14608 27285
rect 15936 27276 15988 27328
rect 16120 27276 16172 27328
rect 16488 27319 16540 27328
rect 16488 27285 16497 27319
rect 16497 27285 16531 27319
rect 16531 27285 16540 27319
rect 16488 27276 16540 27285
rect 16580 27276 16632 27328
rect 18604 27276 18656 27328
rect 18696 27319 18748 27328
rect 18696 27285 18705 27319
rect 18705 27285 18739 27319
rect 18739 27285 18748 27319
rect 18696 27276 18748 27285
rect 21088 27319 21140 27328
rect 21088 27285 21097 27319
rect 21097 27285 21131 27319
rect 21131 27285 21140 27319
rect 21088 27276 21140 27285
rect 24216 27319 24268 27328
rect 24216 27285 24225 27319
rect 24225 27285 24259 27319
rect 24259 27285 24268 27319
rect 24216 27276 24268 27285
rect 24400 27319 24452 27328
rect 24400 27285 24409 27319
rect 24409 27285 24443 27319
rect 24443 27285 24452 27319
rect 24400 27276 24452 27285
rect 27252 27276 27304 27328
rect 27528 27319 27580 27328
rect 27528 27285 27537 27319
rect 27537 27285 27571 27319
rect 27571 27285 27580 27319
rect 27528 27276 27580 27285
rect 4922 27174 4974 27226
rect 4986 27174 5038 27226
rect 5050 27174 5102 27226
rect 5114 27174 5166 27226
rect 5178 27174 5230 27226
rect 5242 27174 5294 27226
rect 10922 27174 10974 27226
rect 10986 27174 11038 27226
rect 11050 27174 11102 27226
rect 11114 27174 11166 27226
rect 11178 27174 11230 27226
rect 11242 27174 11294 27226
rect 16922 27174 16974 27226
rect 16986 27174 17038 27226
rect 17050 27174 17102 27226
rect 17114 27174 17166 27226
rect 17178 27174 17230 27226
rect 17242 27174 17294 27226
rect 22922 27174 22974 27226
rect 22986 27174 23038 27226
rect 23050 27174 23102 27226
rect 23114 27174 23166 27226
rect 23178 27174 23230 27226
rect 23242 27174 23294 27226
rect 28922 27174 28974 27226
rect 28986 27174 29038 27226
rect 29050 27174 29102 27226
rect 29114 27174 29166 27226
rect 29178 27174 29230 27226
rect 29242 27174 29294 27226
rect 9312 27072 9364 27124
rect 10508 27072 10560 27124
rect 15016 27115 15068 27124
rect 15016 27081 15025 27115
rect 15025 27081 15059 27115
rect 15059 27081 15068 27115
rect 15016 27072 15068 27081
rect 17040 27115 17092 27124
rect 17040 27081 17049 27115
rect 17049 27081 17083 27115
rect 17083 27081 17092 27115
rect 17040 27072 17092 27081
rect 18052 27072 18104 27124
rect 18144 27072 18196 27124
rect 18696 27072 18748 27124
rect 21088 27072 21140 27124
rect 23388 27072 23440 27124
rect 24400 27072 24452 27124
rect 26608 27072 26660 27124
rect 27528 27072 27580 27124
rect 11336 27004 11388 27056
rect 6092 26936 6144 26988
rect 8392 26868 8444 26920
rect 13636 26936 13688 26988
rect 14832 27004 14884 27056
rect 15844 27004 15896 27056
rect 15936 27004 15988 27056
rect 16764 27004 16816 27056
rect 9680 26868 9732 26920
rect 10600 26868 10652 26920
rect 12532 26911 12584 26920
rect 12532 26877 12541 26911
rect 12541 26877 12575 26911
rect 12575 26877 12584 26911
rect 12532 26868 12584 26877
rect 13452 26868 13504 26920
rect 14924 26936 14976 26988
rect 15016 26936 15068 26988
rect 16120 26979 16172 26988
rect 16120 26945 16129 26979
rect 16129 26945 16163 26979
rect 16163 26945 16172 26979
rect 16120 26936 16172 26945
rect 16580 26936 16632 26988
rect 17408 27004 17460 27056
rect 17132 26936 17184 26988
rect 18236 27004 18288 27056
rect 17684 26979 17736 26988
rect 17684 26945 17693 26979
rect 17693 26945 17727 26979
rect 17727 26945 17736 26979
rect 17684 26936 17736 26945
rect 17776 26979 17828 26988
rect 17776 26945 17810 26979
rect 17810 26945 17828 26979
rect 17776 26936 17828 26945
rect 18328 26936 18380 26988
rect 20536 26979 20588 26988
rect 20536 26945 20545 26979
rect 20545 26945 20579 26979
rect 20579 26945 20588 26979
rect 20536 26936 20588 26945
rect 23756 26979 23808 26988
rect 23756 26945 23765 26979
rect 23765 26945 23799 26979
rect 23799 26945 23808 26979
rect 23756 26936 23808 26945
rect 29368 27072 29420 27124
rect 28724 26979 28776 26988
rect 28724 26945 28733 26979
rect 28733 26945 28767 26979
rect 28767 26945 28776 26979
rect 28724 26936 28776 26945
rect 14740 26911 14792 26920
rect 14740 26877 14776 26911
rect 14776 26877 14792 26911
rect 14740 26868 14792 26877
rect 12808 26843 12860 26852
rect 12808 26809 12817 26843
rect 12817 26809 12851 26843
rect 12851 26809 12860 26843
rect 12808 26800 12860 26809
rect 15108 26911 15160 26920
rect 15108 26877 15117 26911
rect 15117 26877 15151 26911
rect 15151 26877 15160 26911
rect 15108 26868 15160 26877
rect 16028 26868 16080 26920
rect 6736 26775 6788 26784
rect 6736 26741 6745 26775
rect 6745 26741 6779 26775
rect 6779 26741 6788 26775
rect 6736 26732 6788 26741
rect 15016 26732 15068 26784
rect 15384 26775 15436 26784
rect 15384 26741 15393 26775
rect 15393 26741 15427 26775
rect 15427 26741 15436 26775
rect 15384 26732 15436 26741
rect 16396 26800 16448 26852
rect 16856 26800 16908 26852
rect 18420 26868 18472 26920
rect 19156 26868 19208 26920
rect 20444 26911 20496 26920
rect 20444 26877 20453 26911
rect 20453 26877 20487 26911
rect 20487 26877 20496 26911
rect 20444 26868 20496 26877
rect 19340 26800 19392 26852
rect 25228 26868 25280 26920
rect 25320 26868 25372 26920
rect 27712 26868 27764 26920
rect 18696 26775 18748 26784
rect 18696 26741 18705 26775
rect 18705 26741 18739 26775
rect 18739 26741 18748 26775
rect 18696 26732 18748 26741
rect 18788 26732 18840 26784
rect 21180 26732 21232 26784
rect 27528 26732 27580 26784
rect 27804 26775 27856 26784
rect 27804 26741 27813 26775
rect 27813 26741 27847 26775
rect 27847 26741 27856 26775
rect 27804 26732 27856 26741
rect 4182 26630 4234 26682
rect 4246 26630 4298 26682
rect 4310 26630 4362 26682
rect 4374 26630 4426 26682
rect 4438 26630 4490 26682
rect 4502 26630 4554 26682
rect 10182 26630 10234 26682
rect 10246 26630 10298 26682
rect 10310 26630 10362 26682
rect 10374 26630 10426 26682
rect 10438 26630 10490 26682
rect 10502 26630 10554 26682
rect 16182 26630 16234 26682
rect 16246 26630 16298 26682
rect 16310 26630 16362 26682
rect 16374 26630 16426 26682
rect 16438 26630 16490 26682
rect 16502 26630 16554 26682
rect 22182 26630 22234 26682
rect 22246 26630 22298 26682
rect 22310 26630 22362 26682
rect 22374 26630 22426 26682
rect 22438 26630 22490 26682
rect 22502 26630 22554 26682
rect 28182 26630 28234 26682
rect 28246 26630 28298 26682
rect 28310 26630 28362 26682
rect 28374 26630 28426 26682
rect 28438 26630 28490 26682
rect 28502 26630 28554 26682
rect 8392 26528 8444 26580
rect 9128 26528 9180 26580
rect 18144 26571 18196 26580
rect 18144 26537 18153 26571
rect 18153 26537 18187 26571
rect 18187 26537 18196 26571
rect 18144 26528 18196 26537
rect 18604 26528 18656 26580
rect 18696 26528 18748 26580
rect 19156 26528 19208 26580
rect 27712 26528 27764 26580
rect 27804 26528 27856 26580
rect 28724 26528 28776 26580
rect 14556 26460 14608 26512
rect 14924 26460 14976 26512
rect 16764 26460 16816 26512
rect 18236 26460 18288 26512
rect 9956 26392 10008 26444
rect 7288 26324 7340 26376
rect 14740 26392 14792 26444
rect 15108 26392 15160 26444
rect 16028 26392 16080 26444
rect 17132 26435 17184 26444
rect 17132 26401 17141 26435
rect 17141 26401 17175 26435
rect 17175 26401 17184 26435
rect 17132 26392 17184 26401
rect 17776 26392 17828 26444
rect 13912 26367 13964 26376
rect 13912 26333 13921 26367
rect 13921 26333 13955 26367
rect 13955 26333 13964 26367
rect 13912 26324 13964 26333
rect 14280 26324 14332 26376
rect 3976 26188 4028 26240
rect 7104 26256 7156 26308
rect 7564 26188 7616 26240
rect 8576 26188 8628 26240
rect 11336 26188 11388 26240
rect 13176 26256 13228 26308
rect 17500 26324 17552 26376
rect 18052 26324 18104 26376
rect 15568 26299 15620 26308
rect 15568 26265 15577 26299
rect 15577 26265 15611 26299
rect 15611 26265 15620 26299
rect 15568 26256 15620 26265
rect 15752 26256 15804 26308
rect 17040 26256 17092 26308
rect 17592 26299 17644 26308
rect 17592 26265 17601 26299
rect 17601 26265 17635 26299
rect 17635 26265 17644 26299
rect 17592 26256 17644 26265
rect 17684 26256 17736 26308
rect 18328 26256 18380 26308
rect 24492 26392 24544 26444
rect 25320 26392 25372 26444
rect 27436 26435 27488 26444
rect 27436 26401 27445 26435
rect 27445 26401 27479 26435
rect 27479 26401 27488 26435
rect 27436 26392 27488 26401
rect 23480 26367 23532 26376
rect 23480 26333 23489 26367
rect 23489 26333 23523 26367
rect 23523 26333 23532 26367
rect 23480 26324 23532 26333
rect 23664 26367 23716 26376
rect 23664 26333 23673 26367
rect 23673 26333 23707 26367
rect 23707 26333 23716 26367
rect 23664 26324 23716 26333
rect 24308 26324 24360 26376
rect 15200 26231 15252 26240
rect 15200 26197 15209 26231
rect 15209 26197 15243 26231
rect 15243 26197 15252 26231
rect 15200 26188 15252 26197
rect 16488 26188 16540 26240
rect 18788 26188 18840 26240
rect 19708 26188 19760 26240
rect 20260 26256 20312 26308
rect 26148 26256 26200 26308
rect 31116 26299 31168 26308
rect 31116 26265 31125 26299
rect 31125 26265 31159 26299
rect 31159 26265 31168 26299
rect 31116 26256 31168 26265
rect 31484 26299 31536 26308
rect 31484 26265 31493 26299
rect 31493 26265 31527 26299
rect 31527 26265 31536 26299
rect 31484 26256 31536 26265
rect 20168 26231 20220 26240
rect 20168 26197 20177 26231
rect 20177 26197 20211 26231
rect 20211 26197 20220 26231
rect 20168 26188 20220 26197
rect 23388 26188 23440 26240
rect 24032 26188 24084 26240
rect 24400 26231 24452 26240
rect 24400 26197 24409 26231
rect 24409 26197 24443 26231
rect 24443 26197 24452 26231
rect 24400 26188 24452 26197
rect 26884 26188 26936 26240
rect 27712 26188 27764 26240
rect 4922 26086 4974 26138
rect 4986 26086 5038 26138
rect 5050 26086 5102 26138
rect 5114 26086 5166 26138
rect 5178 26086 5230 26138
rect 5242 26086 5294 26138
rect 10922 26086 10974 26138
rect 10986 26086 11038 26138
rect 11050 26086 11102 26138
rect 11114 26086 11166 26138
rect 11178 26086 11230 26138
rect 11242 26086 11294 26138
rect 16922 26086 16974 26138
rect 16986 26086 17038 26138
rect 17050 26086 17102 26138
rect 17114 26086 17166 26138
rect 17178 26086 17230 26138
rect 17242 26086 17294 26138
rect 22922 26086 22974 26138
rect 22986 26086 23038 26138
rect 23050 26086 23102 26138
rect 23114 26086 23166 26138
rect 23178 26086 23230 26138
rect 23242 26086 23294 26138
rect 28922 26086 28974 26138
rect 28986 26086 29038 26138
rect 29050 26086 29102 26138
rect 29114 26086 29166 26138
rect 29178 26086 29230 26138
rect 29242 26086 29294 26138
rect 6736 26027 6788 26036
rect 6736 25993 6745 26027
rect 6745 25993 6779 26027
rect 6779 25993 6788 26027
rect 6736 25984 6788 25993
rect 7104 25984 7156 26036
rect 7564 26027 7616 26036
rect 7564 25993 7573 26027
rect 7573 25993 7607 26027
rect 7607 25993 7616 26027
rect 7564 25984 7616 25993
rect 5908 25916 5960 25968
rect 8576 25984 8628 26036
rect 13912 25984 13964 26036
rect 14832 25984 14884 26036
rect 14924 25984 14976 26036
rect 16672 25984 16724 26036
rect 18052 25984 18104 26036
rect 21180 25984 21232 26036
rect 22008 25984 22060 26036
rect 25596 25984 25648 26036
rect 15200 25916 15252 25968
rect 15384 25959 15436 25968
rect 15384 25925 15393 25959
rect 15393 25925 15427 25959
rect 15427 25925 15436 25959
rect 15384 25916 15436 25925
rect 19340 25916 19392 25968
rect 4804 25823 4856 25832
rect 4804 25789 4813 25823
rect 4813 25789 4847 25823
rect 4847 25789 4856 25823
rect 4804 25780 4856 25789
rect 6000 25823 6052 25832
rect 6000 25789 6009 25823
rect 6009 25789 6043 25823
rect 6043 25789 6052 25823
rect 6000 25780 6052 25789
rect 9680 25891 9732 25900
rect 9680 25857 9689 25891
rect 9689 25857 9723 25891
rect 9723 25857 9732 25891
rect 9680 25848 9732 25857
rect 9864 25891 9916 25900
rect 9864 25857 9871 25891
rect 9871 25857 9916 25891
rect 9864 25848 9916 25857
rect 10048 25891 10100 25900
rect 10048 25857 10057 25891
rect 10057 25857 10091 25891
rect 10091 25857 10100 25891
rect 10048 25848 10100 25857
rect 10140 25891 10192 25900
rect 10140 25857 10154 25891
rect 10154 25857 10188 25891
rect 10188 25857 10192 25891
rect 10140 25848 10192 25857
rect 10692 25848 10744 25900
rect 14648 25848 14700 25900
rect 18236 25848 18288 25900
rect 22836 25848 22888 25900
rect 5448 25712 5500 25764
rect 8300 25823 8352 25832
rect 8300 25789 8309 25823
rect 8309 25789 8343 25823
rect 8343 25789 8352 25823
rect 8300 25780 8352 25789
rect 13176 25780 13228 25832
rect 14372 25780 14424 25832
rect 22652 25780 22704 25832
rect 23204 25891 23256 25900
rect 23204 25857 23238 25891
rect 23238 25857 23256 25891
rect 23204 25848 23256 25857
rect 25320 25916 25372 25968
rect 24032 25780 24084 25832
rect 29000 25916 29052 25968
rect 29368 25916 29420 25968
rect 4620 25644 4672 25696
rect 5540 25644 5592 25696
rect 11336 25712 11388 25764
rect 11612 25712 11664 25764
rect 24308 25755 24360 25764
rect 24308 25721 24317 25755
rect 24317 25721 24351 25755
rect 24351 25721 24360 25755
rect 24308 25712 24360 25721
rect 9496 25644 9548 25696
rect 10140 25644 10192 25696
rect 11428 25644 11480 25696
rect 12164 25644 12216 25696
rect 15660 25687 15712 25696
rect 15660 25653 15669 25687
rect 15669 25653 15703 25687
rect 15703 25653 15712 25687
rect 15660 25644 15712 25653
rect 25596 25712 25648 25764
rect 26792 25780 26844 25832
rect 26884 25780 26936 25832
rect 25504 25644 25556 25696
rect 25780 25687 25832 25696
rect 25780 25653 25789 25687
rect 25789 25653 25823 25687
rect 25823 25653 25832 25687
rect 25780 25644 25832 25653
rect 26056 25687 26108 25696
rect 26056 25653 26065 25687
rect 26065 25653 26099 25687
rect 26099 25653 26108 25687
rect 26056 25644 26108 25653
rect 27712 25712 27764 25764
rect 29368 25755 29420 25764
rect 29368 25721 29377 25755
rect 29377 25721 29411 25755
rect 29411 25721 29420 25755
rect 29368 25712 29420 25721
rect 26792 25644 26844 25696
rect 4182 25542 4234 25594
rect 4246 25542 4298 25594
rect 4310 25542 4362 25594
rect 4374 25542 4426 25594
rect 4438 25542 4490 25594
rect 4502 25542 4554 25594
rect 10182 25542 10234 25594
rect 10246 25542 10298 25594
rect 10310 25542 10362 25594
rect 10374 25542 10426 25594
rect 10438 25542 10490 25594
rect 10502 25542 10554 25594
rect 16182 25542 16234 25594
rect 16246 25542 16298 25594
rect 16310 25542 16362 25594
rect 16374 25542 16426 25594
rect 16438 25542 16490 25594
rect 16502 25542 16554 25594
rect 22182 25542 22234 25594
rect 22246 25542 22298 25594
rect 22310 25542 22362 25594
rect 22374 25542 22426 25594
rect 22438 25542 22490 25594
rect 22502 25542 22554 25594
rect 28182 25542 28234 25594
rect 28246 25542 28298 25594
rect 28310 25542 28362 25594
rect 28374 25542 28426 25594
rect 28438 25542 28490 25594
rect 28502 25542 28554 25594
rect 5448 25483 5500 25492
rect 5448 25449 5457 25483
rect 5457 25449 5491 25483
rect 5491 25449 5500 25483
rect 5448 25440 5500 25449
rect 6000 25440 6052 25492
rect 5632 25372 5684 25424
rect 3976 25347 4028 25356
rect 3976 25313 3985 25347
rect 3985 25313 4019 25347
rect 4019 25313 4028 25347
rect 3976 25304 4028 25313
rect 5908 25347 5960 25356
rect 5908 25313 5917 25347
rect 5917 25313 5951 25347
rect 5951 25313 5960 25347
rect 5908 25304 5960 25313
rect 6000 25347 6052 25356
rect 6000 25313 6009 25347
rect 6009 25313 6043 25347
rect 6043 25313 6052 25347
rect 6000 25304 6052 25313
rect 9220 25440 9272 25492
rect 9680 25483 9732 25492
rect 9680 25449 9689 25483
rect 9689 25449 9723 25483
rect 9723 25449 9732 25483
rect 9680 25440 9732 25449
rect 20168 25440 20220 25492
rect 8392 25372 8444 25424
rect 9864 25372 9916 25424
rect 10692 25372 10744 25424
rect 6920 25279 6972 25288
rect 6920 25245 6929 25279
rect 6929 25245 6963 25279
rect 6963 25245 6972 25279
rect 6920 25236 6972 25245
rect 7288 25279 7340 25288
rect 7288 25245 7297 25279
rect 7297 25245 7331 25279
rect 7331 25245 7340 25279
rect 7288 25236 7340 25245
rect 8668 25236 8720 25288
rect 4804 25168 4856 25220
rect 7748 25168 7800 25220
rect 8576 25100 8628 25152
rect 8944 25143 8996 25152
rect 8944 25109 8953 25143
rect 8953 25109 8987 25143
rect 8987 25109 8996 25143
rect 8944 25100 8996 25109
rect 9312 25100 9364 25152
rect 9956 25279 10008 25288
rect 9956 25245 9965 25279
rect 9965 25245 9999 25279
rect 9999 25245 10008 25279
rect 9956 25236 10008 25245
rect 12072 25304 12124 25356
rect 22652 25440 22704 25492
rect 23480 25483 23532 25492
rect 23480 25449 23489 25483
rect 23489 25449 23523 25483
rect 23523 25449 23532 25483
rect 23480 25440 23532 25449
rect 23664 25440 23716 25492
rect 26056 25440 26108 25492
rect 24032 25347 24084 25356
rect 24032 25313 24041 25347
rect 24041 25313 24075 25347
rect 24075 25313 24084 25347
rect 24032 25304 24084 25313
rect 24492 25304 24544 25356
rect 25136 25304 25188 25356
rect 10784 25279 10836 25288
rect 10784 25245 10793 25279
rect 10793 25245 10827 25279
rect 10827 25245 10836 25279
rect 10784 25236 10836 25245
rect 18512 25236 18564 25288
rect 19340 25236 19392 25288
rect 19892 25236 19944 25288
rect 24400 25236 24452 25288
rect 10048 25211 10100 25220
rect 10048 25177 10057 25211
rect 10057 25177 10091 25211
rect 10091 25177 10100 25211
rect 10048 25168 10100 25177
rect 11336 25168 11388 25220
rect 16488 25168 16540 25220
rect 25780 25304 25832 25356
rect 9772 25100 9824 25152
rect 10600 25100 10652 25152
rect 12256 25143 12308 25152
rect 12256 25109 12265 25143
rect 12265 25109 12299 25143
rect 12299 25109 12308 25143
rect 12256 25100 12308 25109
rect 19432 25100 19484 25152
rect 21548 25100 21600 25152
rect 29736 25168 29788 25220
rect 25504 25100 25556 25152
rect 26148 25100 26200 25152
rect 4922 24998 4974 25050
rect 4986 24998 5038 25050
rect 5050 24998 5102 25050
rect 5114 24998 5166 25050
rect 5178 24998 5230 25050
rect 5242 24998 5294 25050
rect 10922 24998 10974 25050
rect 10986 24998 11038 25050
rect 11050 24998 11102 25050
rect 11114 24998 11166 25050
rect 11178 24998 11230 25050
rect 11242 24998 11294 25050
rect 16922 24998 16974 25050
rect 16986 24998 17038 25050
rect 17050 24998 17102 25050
rect 17114 24998 17166 25050
rect 17178 24998 17230 25050
rect 17242 24998 17294 25050
rect 22922 24998 22974 25050
rect 22986 24998 23038 25050
rect 23050 24998 23102 25050
rect 23114 24998 23166 25050
rect 23178 24998 23230 25050
rect 23242 24998 23294 25050
rect 28922 24998 28974 25050
rect 28986 24998 29038 25050
rect 29050 24998 29102 25050
rect 29114 24998 29166 25050
rect 29178 24998 29230 25050
rect 29242 24998 29294 25050
rect 4804 24896 4856 24948
rect 5540 24896 5592 24948
rect 7748 24939 7800 24948
rect 7748 24905 7757 24939
rect 7757 24905 7791 24939
rect 7791 24905 7800 24939
rect 7748 24896 7800 24905
rect 8944 24896 8996 24948
rect 11336 24896 11388 24948
rect 12256 24896 12308 24948
rect 4620 24828 4672 24880
rect 3976 24760 4028 24812
rect 940 24692 992 24744
rect 3792 24692 3844 24744
rect 6920 24624 6972 24676
rect 8300 24692 8352 24744
rect 8852 24760 8904 24812
rect 8668 24692 8720 24744
rect 9220 24735 9272 24744
rect 9220 24701 9229 24735
rect 9229 24701 9263 24735
rect 9263 24701 9272 24735
rect 9220 24692 9272 24701
rect 10600 24624 10652 24676
rect 10692 24667 10744 24676
rect 10692 24633 10701 24667
rect 10701 24633 10735 24667
rect 10735 24633 10744 24667
rect 10692 24624 10744 24633
rect 16488 24896 16540 24948
rect 19892 24939 19944 24948
rect 19892 24905 19901 24939
rect 19901 24905 19935 24939
rect 19935 24905 19944 24939
rect 19892 24896 19944 24905
rect 19432 24828 19484 24880
rect 24308 24828 24360 24880
rect 9680 24556 9732 24608
rect 14832 24760 14884 24812
rect 20076 24803 20128 24812
rect 20076 24769 20085 24803
rect 20085 24769 20119 24803
rect 20119 24769 20128 24803
rect 20076 24760 20128 24769
rect 24216 24803 24268 24812
rect 24216 24769 24225 24803
rect 24225 24769 24259 24803
rect 24259 24769 24268 24803
rect 24216 24760 24268 24769
rect 25780 24896 25832 24948
rect 29368 24896 29420 24948
rect 28816 24828 28868 24880
rect 29460 24828 29512 24880
rect 12164 24735 12216 24744
rect 12164 24701 12173 24735
rect 12173 24701 12207 24735
rect 12207 24701 12216 24735
rect 12164 24692 12216 24701
rect 13820 24692 13872 24744
rect 17960 24692 18012 24744
rect 18420 24735 18472 24744
rect 18420 24701 18429 24735
rect 18429 24701 18463 24735
rect 18463 24701 18472 24735
rect 18420 24692 18472 24701
rect 24124 24692 24176 24744
rect 14004 24624 14056 24676
rect 24308 24624 24360 24676
rect 26516 24760 26568 24812
rect 27160 24803 27212 24812
rect 27160 24769 27169 24803
rect 27169 24769 27203 24803
rect 27203 24769 27212 24803
rect 27160 24760 27212 24769
rect 27252 24803 27304 24812
rect 27252 24769 27261 24803
rect 27261 24769 27295 24803
rect 27295 24769 27304 24803
rect 27252 24760 27304 24769
rect 27344 24803 27396 24812
rect 27344 24769 27353 24803
rect 27353 24769 27387 24803
rect 27387 24769 27396 24803
rect 27344 24760 27396 24769
rect 27528 24803 27580 24812
rect 27528 24769 27537 24803
rect 27537 24769 27571 24803
rect 27571 24769 27580 24803
rect 27528 24760 27580 24769
rect 29368 24760 29420 24812
rect 26884 24692 26936 24744
rect 28724 24692 28776 24744
rect 29736 24735 29788 24744
rect 29736 24701 29745 24735
rect 29745 24701 29779 24735
rect 29779 24701 29788 24735
rect 29736 24692 29788 24701
rect 26700 24624 26752 24676
rect 12164 24556 12216 24608
rect 14096 24556 14148 24608
rect 19432 24556 19484 24608
rect 24768 24599 24820 24608
rect 24768 24565 24777 24599
rect 24777 24565 24811 24599
rect 24811 24565 24820 24599
rect 24768 24556 24820 24565
rect 25964 24599 26016 24608
rect 25964 24565 25973 24599
rect 25973 24565 26007 24599
rect 26007 24565 26016 24599
rect 25964 24556 26016 24565
rect 26976 24599 27028 24608
rect 26976 24565 26985 24599
rect 26985 24565 27019 24599
rect 27019 24565 27028 24599
rect 26976 24556 27028 24565
rect 29000 24556 29052 24608
rect 29184 24599 29236 24608
rect 29184 24565 29193 24599
rect 29193 24565 29227 24599
rect 29227 24565 29236 24599
rect 29184 24556 29236 24565
rect 30196 24599 30248 24608
rect 30196 24565 30205 24599
rect 30205 24565 30239 24599
rect 30239 24565 30248 24599
rect 30196 24556 30248 24565
rect 30840 24556 30892 24608
rect 4182 24454 4234 24506
rect 4246 24454 4298 24506
rect 4310 24454 4362 24506
rect 4374 24454 4426 24506
rect 4438 24454 4490 24506
rect 4502 24454 4554 24506
rect 10182 24454 10234 24506
rect 10246 24454 10298 24506
rect 10310 24454 10362 24506
rect 10374 24454 10426 24506
rect 10438 24454 10490 24506
rect 10502 24454 10554 24506
rect 16182 24454 16234 24506
rect 16246 24454 16298 24506
rect 16310 24454 16362 24506
rect 16374 24454 16426 24506
rect 16438 24454 16490 24506
rect 16502 24454 16554 24506
rect 22182 24454 22234 24506
rect 22246 24454 22298 24506
rect 22310 24454 22362 24506
rect 22374 24454 22426 24506
rect 22438 24454 22490 24506
rect 22502 24454 22554 24506
rect 28182 24454 28234 24506
rect 28246 24454 28298 24506
rect 28310 24454 28362 24506
rect 28374 24454 28426 24506
rect 28438 24454 28490 24506
rect 28502 24454 28554 24506
rect 9220 24352 9272 24404
rect 9496 24352 9548 24404
rect 12164 24352 12216 24404
rect 12348 24352 12400 24404
rect 15660 24352 15712 24404
rect 18420 24352 18472 24404
rect 18880 24395 18932 24404
rect 18880 24361 18889 24395
rect 18889 24361 18923 24395
rect 18923 24361 18932 24395
rect 18880 24352 18932 24361
rect 20076 24395 20128 24404
rect 20076 24361 20085 24395
rect 20085 24361 20119 24395
rect 20119 24361 20128 24395
rect 20076 24352 20128 24361
rect 25964 24395 26016 24404
rect 25964 24361 25973 24395
rect 25973 24361 26007 24395
rect 26007 24361 26016 24395
rect 25964 24352 26016 24361
rect 26976 24352 27028 24404
rect 29184 24352 29236 24404
rect 29368 24395 29420 24404
rect 29368 24361 29377 24395
rect 29377 24361 29411 24395
rect 29411 24361 29420 24395
rect 29368 24352 29420 24361
rect 5632 24148 5684 24200
rect 5908 24191 5960 24200
rect 5908 24157 5917 24191
rect 5917 24157 5951 24191
rect 5951 24157 5960 24191
rect 5908 24148 5960 24157
rect 5724 24123 5776 24132
rect 5724 24089 5733 24123
rect 5733 24089 5767 24123
rect 5767 24089 5776 24123
rect 5724 24080 5776 24089
rect 6920 24080 6972 24132
rect 8576 24080 8628 24132
rect 8024 24012 8076 24064
rect 10692 24148 10744 24200
rect 11428 24148 11480 24200
rect 12992 24148 13044 24200
rect 14004 24216 14056 24268
rect 16304 24259 16356 24268
rect 16304 24225 16313 24259
rect 16313 24225 16347 24259
rect 16347 24225 16356 24259
rect 16304 24216 16356 24225
rect 19616 24216 19668 24268
rect 20536 24259 20588 24268
rect 20536 24225 20545 24259
rect 20545 24225 20579 24259
rect 20579 24225 20588 24259
rect 20536 24216 20588 24225
rect 21180 24216 21232 24268
rect 24768 24216 24820 24268
rect 14096 24148 14148 24200
rect 14740 24148 14792 24200
rect 12072 24080 12124 24132
rect 12164 24123 12216 24132
rect 12164 24089 12173 24123
rect 12173 24089 12207 24123
rect 12207 24089 12216 24123
rect 12164 24080 12216 24089
rect 9956 24012 10008 24064
rect 10692 24012 10744 24064
rect 12716 24012 12768 24064
rect 13544 24055 13596 24064
rect 13544 24021 13553 24055
rect 13553 24021 13587 24055
rect 13587 24021 13596 24055
rect 13544 24012 13596 24021
rect 13636 24055 13688 24064
rect 13636 24021 13645 24055
rect 13645 24021 13679 24055
rect 13679 24021 13688 24055
rect 13636 24012 13688 24021
rect 19064 24148 19116 24200
rect 19524 24148 19576 24200
rect 20076 24148 20128 24200
rect 20352 24191 20404 24200
rect 20352 24157 20361 24191
rect 20361 24157 20395 24191
rect 20395 24157 20404 24191
rect 20352 24148 20404 24157
rect 20444 24191 20496 24200
rect 20444 24157 20453 24191
rect 20453 24157 20487 24191
rect 20487 24157 20496 24191
rect 20444 24148 20496 24157
rect 21456 24191 21508 24200
rect 21456 24157 21465 24191
rect 21465 24157 21499 24191
rect 21499 24157 21508 24191
rect 21456 24148 21508 24157
rect 21548 24191 21600 24200
rect 21548 24157 21557 24191
rect 21557 24157 21591 24191
rect 21591 24157 21600 24191
rect 21548 24148 21600 24157
rect 13912 24012 13964 24064
rect 14280 24055 14332 24064
rect 14280 24021 14289 24055
rect 14289 24021 14323 24055
rect 14323 24021 14332 24055
rect 14280 24012 14332 24021
rect 14464 24012 14516 24064
rect 15292 24012 15344 24064
rect 19708 24055 19760 24064
rect 19708 24021 19717 24055
rect 19717 24021 19751 24055
rect 19751 24021 19760 24055
rect 19708 24012 19760 24021
rect 19984 24012 20036 24064
rect 20720 24123 20772 24132
rect 20720 24089 20729 24123
rect 20729 24089 20763 24123
rect 20763 24089 20772 24123
rect 20720 24080 20772 24089
rect 23388 24148 23440 24200
rect 26056 24191 26108 24200
rect 26056 24157 26065 24191
rect 26065 24157 26099 24191
rect 26099 24157 26108 24191
rect 26056 24148 26108 24157
rect 28816 24259 28868 24268
rect 28816 24225 28825 24259
rect 28825 24225 28859 24259
rect 28859 24225 28868 24259
rect 28816 24216 28868 24225
rect 29276 24216 29328 24268
rect 28816 24080 28868 24132
rect 29000 24123 29052 24132
rect 29000 24089 29009 24123
rect 29009 24089 29043 24123
rect 29043 24089 29052 24123
rect 29000 24080 29052 24089
rect 26516 24012 26568 24064
rect 29552 24012 29604 24064
rect 30840 24012 30892 24064
rect 4922 23910 4974 23962
rect 4986 23910 5038 23962
rect 5050 23910 5102 23962
rect 5114 23910 5166 23962
rect 5178 23910 5230 23962
rect 5242 23910 5294 23962
rect 10922 23910 10974 23962
rect 10986 23910 11038 23962
rect 11050 23910 11102 23962
rect 11114 23910 11166 23962
rect 11178 23910 11230 23962
rect 11242 23910 11294 23962
rect 16922 23910 16974 23962
rect 16986 23910 17038 23962
rect 17050 23910 17102 23962
rect 17114 23910 17166 23962
rect 17178 23910 17230 23962
rect 17242 23910 17294 23962
rect 22922 23910 22974 23962
rect 22986 23910 23038 23962
rect 23050 23910 23102 23962
rect 23114 23910 23166 23962
rect 23178 23910 23230 23962
rect 23242 23910 23294 23962
rect 28922 23910 28974 23962
rect 28986 23910 29038 23962
rect 29050 23910 29102 23962
rect 29114 23910 29166 23962
rect 29178 23910 29230 23962
rect 29242 23910 29294 23962
rect 3792 23808 3844 23860
rect 12532 23808 12584 23860
rect 13452 23808 13504 23860
rect 9772 23740 9824 23792
rect 10048 23740 10100 23792
rect 14372 23808 14424 23860
rect 14648 23740 14700 23792
rect 14832 23740 14884 23792
rect 16028 23808 16080 23860
rect 16304 23808 16356 23860
rect 20352 23808 20404 23860
rect 20720 23808 20772 23860
rect 20996 23808 21048 23860
rect 24308 23808 24360 23860
rect 26056 23808 26108 23860
rect 28816 23808 28868 23860
rect 8116 23672 8168 23724
rect 8852 23604 8904 23656
rect 9588 23604 9640 23656
rect 12348 23604 12400 23656
rect 12992 23604 13044 23656
rect 13912 23672 13964 23724
rect 13544 23604 13596 23656
rect 13820 23604 13872 23656
rect 14096 23647 14148 23656
rect 14096 23613 14105 23647
rect 14105 23613 14139 23647
rect 14139 23613 14148 23647
rect 14096 23604 14148 23613
rect 14740 23672 14792 23724
rect 19616 23783 19668 23792
rect 19616 23749 19625 23783
rect 19625 23749 19659 23783
rect 19659 23749 19668 23783
rect 19616 23740 19668 23749
rect 19708 23740 19760 23792
rect 15292 23715 15344 23724
rect 15292 23681 15301 23715
rect 15301 23681 15335 23715
rect 15335 23681 15344 23715
rect 15292 23672 15344 23681
rect 14832 23604 14884 23656
rect 19892 23672 19944 23724
rect 20444 23740 20496 23792
rect 20352 23672 20404 23724
rect 9864 23468 9916 23520
rect 10048 23468 10100 23520
rect 15016 23468 15068 23520
rect 19708 23647 19760 23656
rect 19708 23613 19717 23647
rect 19717 23613 19751 23647
rect 19751 23613 19760 23647
rect 19708 23604 19760 23613
rect 20996 23604 21048 23656
rect 21180 23715 21232 23724
rect 21180 23681 21189 23715
rect 21189 23681 21223 23715
rect 21223 23681 21232 23715
rect 21180 23672 21232 23681
rect 27620 23740 27672 23792
rect 26424 23715 26476 23724
rect 26424 23681 26433 23715
rect 26433 23681 26467 23715
rect 26467 23681 26476 23715
rect 26424 23672 26476 23681
rect 28080 23672 28132 23724
rect 21456 23604 21508 23656
rect 21640 23647 21692 23656
rect 21640 23613 21649 23647
rect 21649 23613 21683 23647
rect 21683 23613 21692 23647
rect 21640 23604 21692 23613
rect 23572 23604 23624 23656
rect 27712 23604 27764 23656
rect 18236 23536 18288 23588
rect 18880 23536 18932 23588
rect 19524 23536 19576 23588
rect 21088 23536 21140 23588
rect 26700 23536 26752 23588
rect 15476 23511 15528 23520
rect 15476 23477 15485 23511
rect 15485 23477 15519 23511
rect 15519 23477 15528 23511
rect 15476 23468 15528 23477
rect 26240 23511 26292 23520
rect 26240 23477 26249 23511
rect 26249 23477 26283 23511
rect 26283 23477 26292 23511
rect 26240 23468 26292 23477
rect 27436 23511 27488 23520
rect 27436 23477 27445 23511
rect 27445 23477 27479 23511
rect 27479 23477 27488 23511
rect 27436 23468 27488 23477
rect 27988 23468 28040 23520
rect 28724 23715 28776 23724
rect 28724 23681 28733 23715
rect 28733 23681 28767 23715
rect 28767 23681 28776 23715
rect 28724 23672 28776 23681
rect 28816 23715 28868 23724
rect 28816 23681 28825 23715
rect 28825 23681 28859 23715
rect 28859 23681 28868 23715
rect 28816 23672 28868 23681
rect 29368 23672 29420 23724
rect 30288 23715 30340 23724
rect 30288 23681 30306 23715
rect 30306 23681 30340 23715
rect 30288 23672 30340 23681
rect 29552 23604 29604 23656
rect 28724 23468 28776 23520
rect 4182 23366 4234 23418
rect 4246 23366 4298 23418
rect 4310 23366 4362 23418
rect 4374 23366 4426 23418
rect 4438 23366 4490 23418
rect 4502 23366 4554 23418
rect 10182 23366 10234 23418
rect 10246 23366 10298 23418
rect 10310 23366 10362 23418
rect 10374 23366 10426 23418
rect 10438 23366 10490 23418
rect 10502 23366 10554 23418
rect 16182 23366 16234 23418
rect 16246 23366 16298 23418
rect 16310 23366 16362 23418
rect 16374 23366 16426 23418
rect 16438 23366 16490 23418
rect 16502 23366 16554 23418
rect 22182 23366 22234 23418
rect 22246 23366 22298 23418
rect 22310 23366 22362 23418
rect 22374 23366 22426 23418
rect 22438 23366 22490 23418
rect 22502 23366 22554 23418
rect 28182 23366 28234 23418
rect 28246 23366 28298 23418
rect 28310 23366 28362 23418
rect 28374 23366 28426 23418
rect 28438 23366 28490 23418
rect 28502 23366 28554 23418
rect 9404 23264 9456 23316
rect 4712 23060 4764 23112
rect 5724 22992 5776 23044
rect 6276 23035 6328 23044
rect 6276 23001 6285 23035
rect 6285 23001 6319 23035
rect 6319 23001 6328 23035
rect 6276 22992 6328 23001
rect 7932 23060 7984 23112
rect 13912 23196 13964 23248
rect 14740 23196 14792 23248
rect 15936 23196 15988 23248
rect 18420 23264 18472 23316
rect 19432 23264 19484 23316
rect 21548 23264 21600 23316
rect 24124 23264 24176 23316
rect 27712 23264 27764 23316
rect 24860 23196 24912 23248
rect 13820 23128 13872 23180
rect 14832 23128 14884 23180
rect 4068 22924 4120 22976
rect 4804 22924 4856 22976
rect 5448 22924 5500 22976
rect 5908 22924 5960 22976
rect 9864 22992 9916 23044
rect 12992 22992 13044 23044
rect 14372 23060 14424 23112
rect 15016 23060 15068 23112
rect 15476 23103 15528 23112
rect 15476 23069 15485 23103
rect 15485 23069 15519 23103
rect 15519 23069 15528 23103
rect 15476 23060 15528 23069
rect 13636 22992 13688 23044
rect 14096 23035 14148 23044
rect 14096 23001 14105 23035
rect 14105 23001 14139 23035
rect 14139 23001 14148 23035
rect 14096 22992 14148 23001
rect 15568 23035 15620 23044
rect 7748 22924 7800 22976
rect 8944 22967 8996 22976
rect 8944 22933 8953 22967
rect 8953 22933 8987 22967
rect 8987 22933 8996 22967
rect 8944 22924 8996 22933
rect 12808 22924 12860 22976
rect 15568 23001 15577 23035
rect 15577 23001 15611 23035
rect 15611 23001 15620 23035
rect 15568 22992 15620 23001
rect 15752 23060 15804 23112
rect 18236 23060 18288 23112
rect 18604 23103 18656 23112
rect 18604 23069 18613 23103
rect 18613 23069 18647 23103
rect 18647 23069 18656 23103
rect 18604 23060 18656 23069
rect 18880 23060 18932 23112
rect 15200 22924 15252 22976
rect 15292 22924 15344 22976
rect 15844 22967 15896 22976
rect 15844 22933 15853 22967
rect 15853 22933 15887 22967
rect 15887 22933 15896 22967
rect 15844 22924 15896 22933
rect 16212 22992 16264 23044
rect 17592 22992 17644 23044
rect 18420 22992 18472 23044
rect 18512 22967 18564 22976
rect 18512 22933 18521 22967
rect 18521 22933 18555 22967
rect 18555 22933 18564 22967
rect 18512 22924 18564 22933
rect 19800 23128 19852 23180
rect 19616 23060 19668 23112
rect 20352 23128 20404 23180
rect 20076 23060 20128 23112
rect 21088 23103 21140 23112
rect 21088 23069 21097 23103
rect 21097 23069 21131 23103
rect 21131 23069 21140 23103
rect 21088 23060 21140 23069
rect 21640 23128 21692 23180
rect 25320 23128 25372 23180
rect 20628 22924 20680 22976
rect 21272 22992 21324 23044
rect 21548 23035 21600 23044
rect 21548 23001 21557 23035
rect 21557 23001 21591 23035
rect 21591 23001 21600 23035
rect 21548 22992 21600 23001
rect 22560 23060 22612 23112
rect 23664 23103 23716 23112
rect 23664 23069 23673 23103
rect 23673 23069 23707 23103
rect 23707 23069 23716 23103
rect 23664 23060 23716 23069
rect 24768 23103 24820 23112
rect 24768 23069 24777 23103
rect 24777 23069 24811 23103
rect 24811 23069 24820 23103
rect 24768 23060 24820 23069
rect 26056 23060 26108 23112
rect 27620 23060 27672 23112
rect 22284 23035 22336 23044
rect 22284 23001 22293 23035
rect 22293 23001 22327 23035
rect 22327 23001 22336 23035
rect 22284 22992 22336 23001
rect 22652 22992 22704 23044
rect 22744 23035 22796 23044
rect 22744 23001 22753 23035
rect 22753 23001 22787 23035
rect 22787 23001 22796 23035
rect 22744 22992 22796 23001
rect 26240 23035 26292 23044
rect 26240 23001 26274 23035
rect 26274 23001 26292 23035
rect 26240 22992 26292 23001
rect 27988 22992 28040 23044
rect 21732 22924 21784 22976
rect 23480 22967 23532 22976
rect 23480 22933 23489 22967
rect 23489 22933 23523 22967
rect 23523 22933 23532 22967
rect 23480 22924 23532 22933
rect 25412 22967 25464 22976
rect 25412 22933 25421 22967
rect 25421 22933 25455 22967
rect 25455 22933 25464 22967
rect 25412 22924 25464 22933
rect 28356 22924 28408 22976
rect 4922 22822 4974 22874
rect 4986 22822 5038 22874
rect 5050 22822 5102 22874
rect 5114 22822 5166 22874
rect 5178 22822 5230 22874
rect 5242 22822 5294 22874
rect 10922 22822 10974 22874
rect 10986 22822 11038 22874
rect 11050 22822 11102 22874
rect 11114 22822 11166 22874
rect 11178 22822 11230 22874
rect 11242 22822 11294 22874
rect 16922 22822 16974 22874
rect 16986 22822 17038 22874
rect 17050 22822 17102 22874
rect 17114 22822 17166 22874
rect 17178 22822 17230 22874
rect 17242 22822 17294 22874
rect 22922 22822 22974 22874
rect 22986 22822 23038 22874
rect 23050 22822 23102 22874
rect 23114 22822 23166 22874
rect 23178 22822 23230 22874
rect 23242 22822 23294 22874
rect 28922 22822 28974 22874
rect 28986 22822 29038 22874
rect 29050 22822 29102 22874
rect 29114 22822 29166 22874
rect 29178 22822 29230 22874
rect 29242 22822 29294 22874
rect 4804 22720 4856 22772
rect 5448 22763 5500 22772
rect 5448 22729 5457 22763
rect 5457 22729 5491 22763
rect 5491 22729 5500 22763
rect 5448 22720 5500 22729
rect 7932 22763 7984 22772
rect 7932 22729 7941 22763
rect 7941 22729 7975 22763
rect 7975 22729 7984 22763
rect 7932 22720 7984 22729
rect 8944 22720 8996 22772
rect 9864 22720 9916 22772
rect 13820 22720 13872 22772
rect 14372 22720 14424 22772
rect 15568 22720 15620 22772
rect 15844 22720 15896 22772
rect 16212 22720 16264 22772
rect 5356 22652 5408 22704
rect 8668 22652 8720 22704
rect 3608 22559 3660 22568
rect 3608 22525 3617 22559
rect 3617 22525 3651 22559
rect 3651 22525 3660 22559
rect 3608 22516 3660 22525
rect 4620 22516 4672 22568
rect 5540 22559 5592 22568
rect 5540 22525 5549 22559
rect 5549 22525 5583 22559
rect 5583 22525 5592 22559
rect 5540 22516 5592 22525
rect 7288 22584 7340 22636
rect 9404 22584 9456 22636
rect 14096 22652 14148 22704
rect 8576 22516 8628 22568
rect 9588 22516 9640 22568
rect 9864 22516 9916 22568
rect 10048 22516 10100 22568
rect 12992 22516 13044 22568
rect 13912 22584 13964 22636
rect 15568 22627 15620 22636
rect 14096 22516 14148 22568
rect 15568 22593 15577 22627
rect 15577 22593 15611 22627
rect 15611 22593 15620 22627
rect 15568 22584 15620 22593
rect 16028 22584 16080 22636
rect 17960 22720 18012 22772
rect 19340 22652 19392 22704
rect 20812 22720 20864 22772
rect 15936 22559 15988 22568
rect 15936 22525 15945 22559
rect 15945 22525 15979 22559
rect 15979 22525 15988 22559
rect 15936 22516 15988 22525
rect 19064 22584 19116 22636
rect 19616 22584 19668 22636
rect 19984 22584 20036 22636
rect 20076 22584 20128 22636
rect 22836 22652 22888 22704
rect 8024 22423 8076 22432
rect 8024 22389 8033 22423
rect 8033 22389 8067 22423
rect 8067 22389 8076 22423
rect 8024 22380 8076 22389
rect 11060 22380 11112 22432
rect 12164 22380 12216 22432
rect 14648 22380 14700 22432
rect 15200 22380 15252 22432
rect 15844 22380 15896 22432
rect 18604 22448 18656 22500
rect 20904 22584 20956 22636
rect 21732 22584 21784 22636
rect 22560 22627 22612 22636
rect 22560 22593 22569 22627
rect 22569 22593 22603 22627
rect 22603 22593 22612 22627
rect 22560 22584 22612 22593
rect 22652 22627 22704 22636
rect 22652 22593 22661 22627
rect 22661 22593 22695 22627
rect 22695 22593 22704 22627
rect 22652 22584 22704 22593
rect 23480 22720 23532 22772
rect 23664 22720 23716 22772
rect 25412 22720 25464 22772
rect 23848 22652 23900 22704
rect 21456 22516 21508 22568
rect 22284 22516 22336 22568
rect 25228 22559 25280 22568
rect 25228 22525 25237 22559
rect 25237 22525 25271 22559
rect 25271 22525 25280 22559
rect 25228 22516 25280 22525
rect 27712 22720 27764 22772
rect 28080 22720 28132 22772
rect 28632 22720 28684 22772
rect 28356 22652 28408 22704
rect 27160 22584 27212 22636
rect 27344 22584 27396 22636
rect 26884 22516 26936 22568
rect 28724 22516 28776 22568
rect 21272 22380 21324 22432
rect 27988 22448 28040 22500
rect 24768 22380 24820 22432
rect 26792 22423 26844 22432
rect 26792 22389 26801 22423
rect 26801 22389 26835 22423
rect 26835 22389 26844 22423
rect 26792 22380 26844 22389
rect 4182 22278 4234 22330
rect 4246 22278 4298 22330
rect 4310 22278 4362 22330
rect 4374 22278 4426 22330
rect 4438 22278 4490 22330
rect 4502 22278 4554 22330
rect 10182 22278 10234 22330
rect 10246 22278 10298 22330
rect 10310 22278 10362 22330
rect 10374 22278 10426 22330
rect 10438 22278 10490 22330
rect 10502 22278 10554 22330
rect 16182 22278 16234 22330
rect 16246 22278 16298 22330
rect 16310 22278 16362 22330
rect 16374 22278 16426 22330
rect 16438 22278 16490 22330
rect 16502 22278 16554 22330
rect 22182 22278 22234 22330
rect 22246 22278 22298 22330
rect 22310 22278 22362 22330
rect 22374 22278 22426 22330
rect 22438 22278 22490 22330
rect 22502 22278 22554 22330
rect 28182 22278 28234 22330
rect 28246 22278 28298 22330
rect 28310 22278 28362 22330
rect 28374 22278 28426 22330
rect 28438 22278 28490 22330
rect 28502 22278 28554 22330
rect 4712 22176 4764 22228
rect 7288 22219 7340 22228
rect 7288 22185 7297 22219
rect 7297 22185 7331 22219
rect 7331 22185 7340 22219
rect 7288 22176 7340 22185
rect 8024 22176 8076 22228
rect 10140 22176 10192 22228
rect 5816 22108 5868 22160
rect 6000 22108 6052 22160
rect 3608 21972 3660 22024
rect 5356 21972 5408 22024
rect 9588 22040 9640 22092
rect 10232 22108 10284 22160
rect 10784 22108 10836 22160
rect 15568 22108 15620 22160
rect 19984 22176 20036 22228
rect 21456 22219 21508 22228
rect 21456 22185 21465 22219
rect 21465 22185 21499 22219
rect 21499 22185 21508 22219
rect 21456 22176 21508 22185
rect 21640 22176 21692 22228
rect 21272 22108 21324 22160
rect 24032 22108 24084 22160
rect 4068 21947 4120 21956
rect 4068 21913 4102 21947
rect 4102 21913 4120 21947
rect 4068 21904 4120 21913
rect 7748 22015 7800 22024
rect 7748 21981 7757 22015
rect 7757 21981 7791 22015
rect 7791 21981 7800 22015
rect 7748 21972 7800 21981
rect 7932 22015 7984 22024
rect 7932 21981 7941 22015
rect 7941 21981 7975 22015
rect 7975 21981 7984 22015
rect 7932 21972 7984 21981
rect 8024 22015 8076 22024
rect 8024 21981 8033 22015
rect 8033 21981 8067 22015
rect 8067 21981 8076 22015
rect 8024 21972 8076 21981
rect 8944 21972 8996 22024
rect 15752 22040 15804 22092
rect 15844 22040 15896 22092
rect 5632 21879 5684 21888
rect 5632 21845 5641 21879
rect 5641 21845 5675 21879
rect 5675 21845 5684 21879
rect 5632 21836 5684 21845
rect 6092 21836 6144 21888
rect 6276 21836 6328 21888
rect 6552 21879 6604 21888
rect 6552 21845 6561 21879
rect 6561 21845 6595 21879
rect 6595 21845 6604 21879
rect 6552 21836 6604 21845
rect 7196 21836 7248 21888
rect 8484 21836 8536 21888
rect 9220 21904 9272 21956
rect 9404 21904 9456 21956
rect 10416 21879 10468 21888
rect 10416 21845 10425 21879
rect 10425 21845 10459 21879
rect 10459 21845 10468 21879
rect 10416 21836 10468 21845
rect 10600 22015 10652 22024
rect 10600 21981 10609 22015
rect 10609 21981 10643 22015
rect 10643 21981 10652 22015
rect 10600 21972 10652 21981
rect 11060 22015 11112 22024
rect 11060 21981 11069 22015
rect 11069 21981 11103 22015
rect 11103 21981 11112 22015
rect 11060 21972 11112 21981
rect 16120 22015 16172 22024
rect 16120 21981 16129 22015
rect 16129 21981 16163 22015
rect 16163 21981 16172 22015
rect 16120 21972 16172 21981
rect 18512 21972 18564 22024
rect 19616 21972 19668 22024
rect 21732 22040 21784 22092
rect 22836 22083 22888 22092
rect 22836 22049 22845 22083
rect 22845 22049 22879 22083
rect 22879 22049 22888 22083
rect 22836 22040 22888 22049
rect 24860 22083 24912 22092
rect 24860 22049 24869 22083
rect 24869 22049 24903 22083
rect 24903 22049 24912 22083
rect 24860 22040 24912 22049
rect 26424 22040 26476 22092
rect 27528 22083 27580 22092
rect 27528 22049 27537 22083
rect 27537 22049 27571 22083
rect 27571 22049 27580 22083
rect 27528 22040 27580 22049
rect 10784 21904 10836 21956
rect 11336 21904 11388 21956
rect 19984 21947 20036 21956
rect 19984 21913 19993 21947
rect 19993 21913 20027 21947
rect 20027 21913 20036 21947
rect 19984 21904 20036 21913
rect 20720 21947 20772 21956
rect 20720 21913 20729 21947
rect 20729 21913 20763 21947
rect 20763 21913 20772 21947
rect 20720 21904 20772 21913
rect 17316 21836 17368 21888
rect 23480 21904 23532 21956
rect 23664 21836 23716 21888
rect 24216 21879 24268 21888
rect 24216 21845 24225 21879
rect 24225 21845 24259 21879
rect 24259 21845 24268 21879
rect 24216 21836 24268 21845
rect 24768 21879 24820 21888
rect 24768 21845 24777 21879
rect 24777 21845 24811 21879
rect 24811 21845 24820 21879
rect 24768 21836 24820 21845
rect 25320 21904 25372 21956
rect 26148 21904 26200 21956
rect 26240 21836 26292 21888
rect 27436 21972 27488 22024
rect 29644 21972 29696 22024
rect 27436 21879 27488 21888
rect 27436 21845 27445 21879
rect 27445 21845 27479 21879
rect 27479 21845 27488 21879
rect 27436 21836 27488 21845
rect 29552 21879 29604 21888
rect 29552 21845 29561 21879
rect 29561 21845 29595 21879
rect 29595 21845 29604 21879
rect 29552 21836 29604 21845
rect 4922 21734 4974 21786
rect 4986 21734 5038 21786
rect 5050 21734 5102 21786
rect 5114 21734 5166 21786
rect 5178 21734 5230 21786
rect 5242 21734 5294 21786
rect 10922 21734 10974 21786
rect 10986 21734 11038 21786
rect 11050 21734 11102 21786
rect 11114 21734 11166 21786
rect 11178 21734 11230 21786
rect 11242 21734 11294 21786
rect 16922 21734 16974 21786
rect 16986 21734 17038 21786
rect 17050 21734 17102 21786
rect 17114 21734 17166 21786
rect 17178 21734 17230 21786
rect 17242 21734 17294 21786
rect 22922 21734 22974 21786
rect 22986 21734 23038 21786
rect 23050 21734 23102 21786
rect 23114 21734 23166 21786
rect 23178 21734 23230 21786
rect 23242 21734 23294 21786
rect 28922 21734 28974 21786
rect 28986 21734 29038 21786
rect 29050 21734 29102 21786
rect 29114 21734 29166 21786
rect 29178 21734 29230 21786
rect 29242 21734 29294 21786
rect 5356 21632 5408 21684
rect 6552 21632 6604 21684
rect 5540 21564 5592 21616
rect 6092 21564 6144 21616
rect 7104 21632 7156 21684
rect 8668 21607 8720 21616
rect 8668 21573 8677 21607
rect 8677 21573 8711 21607
rect 8711 21573 8720 21607
rect 8668 21564 8720 21573
rect 8760 21564 8812 21616
rect 9588 21675 9640 21684
rect 9588 21641 9597 21675
rect 9597 21641 9631 21675
rect 9631 21641 9640 21675
rect 9588 21632 9640 21641
rect 10784 21632 10836 21684
rect 6184 21496 6236 21548
rect 7380 21496 7432 21548
rect 7840 21496 7892 21548
rect 8208 21496 8260 21548
rect 8852 21496 8904 21548
rect 7196 21428 7248 21480
rect 9496 21496 9548 21548
rect 10048 21496 10100 21548
rect 10416 21564 10468 21616
rect 12716 21675 12768 21684
rect 12716 21641 12725 21675
rect 12725 21641 12759 21675
rect 12759 21641 12768 21675
rect 12716 21632 12768 21641
rect 9864 21428 9916 21480
rect 13360 21496 13412 21548
rect 17592 21632 17644 21684
rect 23480 21675 23532 21684
rect 23480 21641 23489 21675
rect 23489 21641 23523 21675
rect 23523 21641 23532 21675
rect 23480 21632 23532 21641
rect 18604 21496 18656 21548
rect 23848 21564 23900 21616
rect 24124 21607 24176 21616
rect 24124 21573 24133 21607
rect 24133 21573 24167 21607
rect 24167 21573 24176 21607
rect 24124 21564 24176 21573
rect 24216 21607 24268 21616
rect 24216 21573 24225 21607
rect 24225 21573 24259 21607
rect 24259 21573 24268 21607
rect 24216 21564 24268 21573
rect 23664 21539 23716 21548
rect 23664 21505 23673 21539
rect 23673 21505 23707 21539
rect 23707 21505 23716 21539
rect 23664 21496 23716 21505
rect 24308 21539 24360 21548
rect 24308 21505 24317 21539
rect 24317 21505 24351 21539
rect 24351 21505 24360 21539
rect 24308 21496 24360 21505
rect 24768 21632 24820 21684
rect 29552 21675 29604 21684
rect 29552 21641 29561 21675
rect 29561 21641 29595 21675
rect 29595 21641 29604 21675
rect 29552 21632 29604 21641
rect 24860 21564 24912 21616
rect 25320 21607 25372 21616
rect 25320 21573 25329 21607
rect 25329 21573 25363 21607
rect 25363 21573 25372 21607
rect 25320 21564 25372 21573
rect 26056 21607 26108 21616
rect 26056 21573 26065 21607
rect 26065 21573 26099 21607
rect 26099 21573 26108 21607
rect 26056 21564 26108 21573
rect 27436 21564 27488 21616
rect 27988 21496 28040 21548
rect 24676 21428 24728 21480
rect 26792 21428 26844 21480
rect 29828 21428 29880 21480
rect 6368 21335 6420 21344
rect 6368 21301 6377 21335
rect 6377 21301 6411 21335
rect 6411 21301 6420 21335
rect 6368 21292 6420 21301
rect 9312 21292 9364 21344
rect 10692 21292 10744 21344
rect 12808 21360 12860 21412
rect 30104 21428 30156 21480
rect 11520 21335 11572 21344
rect 11520 21301 11529 21335
rect 11529 21301 11563 21335
rect 11563 21301 11572 21335
rect 11520 21292 11572 21301
rect 13268 21335 13320 21344
rect 13268 21301 13277 21335
rect 13277 21301 13311 21335
rect 13311 21301 13320 21335
rect 13268 21292 13320 21301
rect 17316 21292 17368 21344
rect 26976 21335 27028 21344
rect 26976 21301 26985 21335
rect 26985 21301 27019 21335
rect 27019 21301 27028 21335
rect 26976 21292 27028 21301
rect 29000 21292 29052 21344
rect 30656 21292 30708 21344
rect 4182 21190 4234 21242
rect 4246 21190 4298 21242
rect 4310 21190 4362 21242
rect 4374 21190 4426 21242
rect 4438 21190 4490 21242
rect 4502 21190 4554 21242
rect 10182 21190 10234 21242
rect 10246 21190 10298 21242
rect 10310 21190 10362 21242
rect 10374 21190 10426 21242
rect 10438 21190 10490 21242
rect 10502 21190 10554 21242
rect 16182 21190 16234 21242
rect 16246 21190 16298 21242
rect 16310 21190 16362 21242
rect 16374 21190 16426 21242
rect 16438 21190 16490 21242
rect 16502 21190 16554 21242
rect 22182 21190 22234 21242
rect 22246 21190 22298 21242
rect 22310 21190 22362 21242
rect 22374 21190 22426 21242
rect 22438 21190 22490 21242
rect 22502 21190 22554 21242
rect 28182 21190 28234 21242
rect 28246 21190 28298 21242
rect 28310 21190 28362 21242
rect 28374 21190 28426 21242
rect 28438 21190 28490 21242
rect 28502 21190 28554 21242
rect 5632 21088 5684 21140
rect 6184 21131 6236 21140
rect 6184 21097 6193 21131
rect 6193 21097 6227 21131
rect 6227 21097 6236 21131
rect 6184 21088 6236 21097
rect 6368 21088 6420 21140
rect 8944 21131 8996 21140
rect 8944 21097 8953 21131
rect 8953 21097 8987 21131
rect 8987 21097 8996 21131
rect 8944 21088 8996 21097
rect 10600 21131 10652 21140
rect 10600 21097 10609 21131
rect 10609 21097 10643 21131
rect 10643 21097 10652 21131
rect 10600 21088 10652 21097
rect 12532 21088 12584 21140
rect 15292 21088 15344 21140
rect 23848 21088 23900 21140
rect 26976 21088 27028 21140
rect 6276 20952 6328 21004
rect 10048 21020 10100 21072
rect 10968 21020 11020 21072
rect 9680 20952 9732 21004
rect 10876 20952 10928 21004
rect 8484 20927 8536 20936
rect 8484 20893 8502 20927
rect 8502 20893 8536 20927
rect 8484 20884 8536 20893
rect 9864 20884 9916 20936
rect 11520 21020 11572 21072
rect 28080 21020 28132 21072
rect 11428 20952 11480 21004
rect 12256 20952 12308 21004
rect 14924 20952 14976 21004
rect 24952 20952 25004 21004
rect 11244 20884 11296 20936
rect 11336 20884 11388 20936
rect 12164 20927 12216 20936
rect 12164 20893 12173 20927
rect 12173 20893 12207 20927
rect 12207 20893 12216 20927
rect 12164 20884 12216 20893
rect 8392 20816 8444 20868
rect 9220 20816 9272 20868
rect 14188 20884 14240 20936
rect 25044 20884 25096 20936
rect 26516 20884 26568 20936
rect 27068 20952 27120 21004
rect 27436 20927 27488 20936
rect 27436 20893 27445 20927
rect 27445 20893 27479 20927
rect 27479 20893 27488 20927
rect 29644 21088 29696 21140
rect 29552 20952 29604 21004
rect 29736 20952 29788 21004
rect 27436 20884 27488 20893
rect 29000 20927 29052 20936
rect 29000 20893 29009 20927
rect 29009 20893 29043 20927
rect 29043 20893 29052 20927
rect 29000 20884 29052 20893
rect 30656 20927 30708 20936
rect 30656 20893 30674 20927
rect 30674 20893 30708 20927
rect 30656 20884 30708 20893
rect 12900 20859 12952 20868
rect 12900 20825 12909 20859
rect 12909 20825 12943 20859
rect 12943 20825 12952 20859
rect 12900 20816 12952 20825
rect 8760 20748 8812 20800
rect 9312 20791 9364 20800
rect 9312 20757 9321 20791
rect 9321 20757 9355 20791
rect 9355 20757 9364 20791
rect 9312 20748 9364 20757
rect 10876 20748 10928 20800
rect 12624 20748 12676 20800
rect 14188 20791 14240 20800
rect 14188 20757 14197 20791
rect 14197 20757 14231 20791
rect 14231 20757 14240 20791
rect 14188 20748 14240 20757
rect 25320 20791 25372 20800
rect 25320 20757 25329 20791
rect 25329 20757 25363 20791
rect 25363 20757 25372 20791
rect 25320 20748 25372 20757
rect 27252 20816 27304 20868
rect 27896 20816 27948 20868
rect 28080 20816 28132 20868
rect 28632 20816 28684 20868
rect 26700 20748 26752 20800
rect 26976 20791 27028 20800
rect 26976 20757 26985 20791
rect 26985 20757 27019 20791
rect 27019 20757 27028 20791
rect 26976 20748 27028 20757
rect 30564 20748 30616 20800
rect 31116 20816 31168 20868
rect 31024 20791 31076 20800
rect 31024 20757 31033 20791
rect 31033 20757 31067 20791
rect 31067 20757 31076 20791
rect 31024 20748 31076 20757
rect 4922 20646 4974 20698
rect 4986 20646 5038 20698
rect 5050 20646 5102 20698
rect 5114 20646 5166 20698
rect 5178 20646 5230 20698
rect 5242 20646 5294 20698
rect 10922 20646 10974 20698
rect 10986 20646 11038 20698
rect 11050 20646 11102 20698
rect 11114 20646 11166 20698
rect 11178 20646 11230 20698
rect 11242 20646 11294 20698
rect 16922 20646 16974 20698
rect 16986 20646 17038 20698
rect 17050 20646 17102 20698
rect 17114 20646 17166 20698
rect 17178 20646 17230 20698
rect 17242 20646 17294 20698
rect 22922 20646 22974 20698
rect 22986 20646 23038 20698
rect 23050 20646 23102 20698
rect 23114 20646 23166 20698
rect 23178 20646 23230 20698
rect 23242 20646 23294 20698
rect 28922 20646 28974 20698
rect 28986 20646 29038 20698
rect 29050 20646 29102 20698
rect 29114 20646 29166 20698
rect 29178 20646 29230 20698
rect 29242 20646 29294 20698
rect 9312 20544 9364 20596
rect 10784 20544 10836 20596
rect 11428 20544 11480 20596
rect 13360 20544 13412 20596
rect 8300 20476 8352 20528
rect 7472 20451 7524 20460
rect 7472 20417 7481 20451
rect 7481 20417 7515 20451
rect 7515 20417 7524 20451
rect 7472 20408 7524 20417
rect 7748 20408 7800 20460
rect 8760 20408 8812 20460
rect 9496 20451 9548 20460
rect 9496 20417 9505 20451
rect 9505 20417 9539 20451
rect 9539 20417 9548 20451
rect 9496 20408 9548 20417
rect 6920 20340 6972 20392
rect 8852 20340 8904 20392
rect 7288 20247 7340 20256
rect 7288 20213 7297 20247
rect 7297 20213 7331 20247
rect 7331 20213 7340 20247
rect 7288 20204 7340 20213
rect 9496 20204 9548 20256
rect 9772 20408 9824 20460
rect 13268 20476 13320 20528
rect 14188 20476 14240 20528
rect 11520 20340 11572 20392
rect 12900 20383 12952 20392
rect 12900 20349 12909 20383
rect 12909 20349 12943 20383
rect 12943 20349 12952 20383
rect 12900 20340 12952 20349
rect 9772 20272 9824 20324
rect 12532 20272 12584 20324
rect 12348 20204 12400 20256
rect 14556 20204 14608 20256
rect 25044 20587 25096 20596
rect 25044 20553 25053 20587
rect 25053 20553 25087 20587
rect 25087 20553 25096 20587
rect 25044 20544 25096 20553
rect 25320 20544 25372 20596
rect 26976 20544 27028 20596
rect 27896 20587 27948 20596
rect 27896 20553 27905 20587
rect 27905 20553 27939 20587
rect 27939 20553 27948 20587
rect 27896 20544 27948 20553
rect 29000 20544 29052 20596
rect 30104 20544 30156 20596
rect 26148 20476 26200 20528
rect 23940 20451 23992 20460
rect 23940 20417 23974 20451
rect 23974 20417 23992 20451
rect 23940 20408 23992 20417
rect 24952 20408 25004 20460
rect 27252 20476 27304 20528
rect 31024 20476 31076 20528
rect 30564 20408 30616 20460
rect 25228 20340 25280 20392
rect 26240 20340 26292 20392
rect 25136 20247 25188 20256
rect 25136 20213 25145 20247
rect 25145 20213 25179 20247
rect 25179 20213 25188 20247
rect 25136 20204 25188 20213
rect 26332 20247 26384 20256
rect 26332 20213 26341 20247
rect 26341 20213 26375 20247
rect 26375 20213 26384 20247
rect 26332 20204 26384 20213
rect 29368 20272 29420 20324
rect 31208 20204 31260 20256
rect 4182 20102 4234 20154
rect 4246 20102 4298 20154
rect 4310 20102 4362 20154
rect 4374 20102 4426 20154
rect 4438 20102 4490 20154
rect 4502 20102 4554 20154
rect 10182 20102 10234 20154
rect 10246 20102 10298 20154
rect 10310 20102 10362 20154
rect 10374 20102 10426 20154
rect 10438 20102 10490 20154
rect 10502 20102 10554 20154
rect 16182 20102 16234 20154
rect 16246 20102 16298 20154
rect 16310 20102 16362 20154
rect 16374 20102 16426 20154
rect 16438 20102 16490 20154
rect 16502 20102 16554 20154
rect 22182 20102 22234 20154
rect 22246 20102 22298 20154
rect 22310 20102 22362 20154
rect 22374 20102 22426 20154
rect 22438 20102 22490 20154
rect 22502 20102 22554 20154
rect 28182 20102 28234 20154
rect 28246 20102 28298 20154
rect 28310 20102 28362 20154
rect 28374 20102 28426 20154
rect 28438 20102 28490 20154
rect 28502 20102 28554 20154
rect 23940 20000 23992 20052
rect 25136 20000 25188 20052
rect 27252 20000 27304 20052
rect 27988 20000 28040 20052
rect 4712 19864 4764 19916
rect 5816 19864 5868 19916
rect 9496 19907 9548 19916
rect 9496 19873 9505 19907
rect 9505 19873 9539 19907
rect 9539 19873 9548 19907
rect 9496 19864 9548 19873
rect 18972 19907 19024 19916
rect 18972 19873 18981 19907
rect 18981 19873 19015 19907
rect 19015 19873 19024 19907
rect 18972 19864 19024 19873
rect 20444 19864 20496 19916
rect 22008 19907 22060 19916
rect 22008 19873 22017 19907
rect 22017 19873 22051 19907
rect 22051 19873 22060 19907
rect 22008 19864 22060 19873
rect 5540 19796 5592 19848
rect 6920 19796 6972 19848
rect 7288 19839 7340 19848
rect 7288 19805 7322 19839
rect 7322 19805 7340 19839
rect 7288 19796 7340 19805
rect 12164 19796 12216 19848
rect 12256 19839 12308 19848
rect 12256 19805 12265 19839
rect 12265 19805 12299 19839
rect 12299 19805 12308 19839
rect 12256 19796 12308 19805
rect 12900 19796 12952 19848
rect 17684 19839 17736 19848
rect 17684 19805 17693 19839
rect 17693 19805 17727 19839
rect 17727 19805 17736 19839
rect 17684 19796 17736 19805
rect 20720 19839 20772 19848
rect 20720 19805 20729 19839
rect 20729 19805 20763 19839
rect 20763 19805 20772 19839
rect 20720 19796 20772 19805
rect 21180 19839 21232 19848
rect 21180 19805 21189 19839
rect 21189 19805 21223 19839
rect 21223 19805 21232 19839
rect 21180 19796 21232 19805
rect 22836 19839 22888 19848
rect 22836 19805 22845 19839
rect 22845 19805 22879 19839
rect 22879 19805 22888 19839
rect 22836 19796 22888 19805
rect 31852 19932 31904 19984
rect 26148 19796 26200 19848
rect 26332 19839 26384 19848
rect 26332 19805 26366 19839
rect 26366 19805 26384 19839
rect 26332 19796 26384 19805
rect 28724 19839 28776 19848
rect 28724 19805 28728 19839
rect 28728 19805 28762 19839
rect 28762 19805 28776 19839
rect 28724 19796 28776 19805
rect 29000 19796 29052 19848
rect 22744 19728 22796 19780
rect 23664 19728 23716 19780
rect 27344 19728 27396 19780
rect 28908 19771 28960 19780
rect 28908 19737 28917 19771
rect 28917 19737 28951 19771
rect 28951 19737 28960 19771
rect 28908 19728 28960 19737
rect 29368 19796 29420 19848
rect 29644 19796 29696 19848
rect 31208 19839 31260 19848
rect 31208 19805 31217 19839
rect 31217 19805 31251 19839
rect 31251 19805 31260 19839
rect 31208 19796 31260 19805
rect 3148 19660 3200 19712
rect 4896 19660 4948 19712
rect 8944 19703 8996 19712
rect 8944 19669 8953 19703
rect 8953 19669 8987 19703
rect 8987 19669 8996 19703
rect 8944 19660 8996 19669
rect 11336 19703 11388 19712
rect 11336 19669 11345 19703
rect 11345 19669 11379 19703
rect 11379 19669 11388 19703
rect 11336 19660 11388 19669
rect 12072 19703 12124 19712
rect 12072 19669 12081 19703
rect 12081 19669 12115 19703
rect 12115 19669 12124 19703
rect 12072 19660 12124 19669
rect 12808 19703 12860 19712
rect 12808 19669 12817 19703
rect 12817 19669 12851 19703
rect 12851 19669 12860 19703
rect 12808 19660 12860 19669
rect 17500 19703 17552 19712
rect 17500 19669 17509 19703
rect 17509 19669 17543 19703
rect 17543 19669 17552 19703
rect 17500 19660 17552 19669
rect 18328 19703 18380 19712
rect 18328 19669 18337 19703
rect 18337 19669 18371 19703
rect 18371 19669 18380 19703
rect 18328 19660 18380 19669
rect 20168 19703 20220 19712
rect 20168 19669 20177 19703
rect 20177 19669 20211 19703
rect 20211 19669 20220 19703
rect 20168 19660 20220 19669
rect 20996 19703 21048 19712
rect 20996 19669 21005 19703
rect 21005 19669 21039 19703
rect 21039 19669 21048 19703
rect 20996 19660 21048 19669
rect 21456 19703 21508 19712
rect 21456 19669 21465 19703
rect 21465 19669 21499 19703
rect 21499 19669 21508 19703
rect 21456 19660 21508 19669
rect 21640 19660 21692 19712
rect 29460 19660 29512 19712
rect 4922 19558 4974 19610
rect 4986 19558 5038 19610
rect 5050 19558 5102 19610
rect 5114 19558 5166 19610
rect 5178 19558 5230 19610
rect 5242 19558 5294 19610
rect 10922 19558 10974 19610
rect 10986 19558 11038 19610
rect 11050 19558 11102 19610
rect 11114 19558 11166 19610
rect 11178 19558 11230 19610
rect 11242 19558 11294 19610
rect 16922 19558 16974 19610
rect 16986 19558 17038 19610
rect 17050 19558 17102 19610
rect 17114 19558 17166 19610
rect 17178 19558 17230 19610
rect 17242 19558 17294 19610
rect 22922 19558 22974 19610
rect 22986 19558 23038 19610
rect 23050 19558 23102 19610
rect 23114 19558 23166 19610
rect 23178 19558 23230 19610
rect 23242 19558 23294 19610
rect 28922 19558 28974 19610
rect 28986 19558 29038 19610
rect 29050 19558 29102 19610
rect 29114 19558 29166 19610
rect 29178 19558 29230 19610
rect 29242 19558 29294 19610
rect 5172 19456 5224 19508
rect 5540 19456 5592 19508
rect 7472 19456 7524 19508
rect 8944 19456 8996 19508
rect 3056 19320 3108 19372
rect 3976 19363 4028 19372
rect 3976 19329 3985 19363
rect 3985 19329 4019 19363
rect 4019 19329 4028 19363
rect 3976 19320 4028 19329
rect 4252 19363 4304 19372
rect 4252 19329 4286 19363
rect 4286 19329 4304 19363
rect 4252 19320 4304 19329
rect 6000 19363 6052 19372
rect 6000 19329 6009 19363
rect 6009 19329 6043 19363
rect 6043 19329 6052 19363
rect 6000 19320 6052 19329
rect 6920 19320 6972 19372
rect 9864 19320 9916 19372
rect 10600 19320 10652 19372
rect 11520 19363 11572 19372
rect 11520 19329 11529 19363
rect 11529 19329 11563 19363
rect 11563 19329 11572 19363
rect 11520 19320 11572 19329
rect 12072 19456 12124 19508
rect 12900 19499 12952 19508
rect 12900 19465 12909 19499
rect 12909 19465 12943 19499
rect 12943 19465 12952 19499
rect 12900 19456 12952 19465
rect 18972 19456 19024 19508
rect 12440 19388 12492 19440
rect 14372 19388 14424 19440
rect 14648 19388 14700 19440
rect 12164 19320 12216 19372
rect 15936 19388 15988 19440
rect 17500 19431 17552 19440
rect 17500 19397 17534 19431
rect 17534 19397 17552 19431
rect 17500 19388 17552 19397
rect 8208 19252 8260 19304
rect 8300 19295 8352 19304
rect 8300 19261 8309 19295
rect 8309 19261 8343 19295
rect 8343 19261 8352 19295
rect 8300 19252 8352 19261
rect 7748 19227 7800 19236
rect 7748 19193 7757 19227
rect 7757 19193 7791 19227
rect 7791 19193 7800 19227
rect 7748 19184 7800 19193
rect 13452 19295 13504 19304
rect 13452 19261 13461 19295
rect 13461 19261 13495 19295
rect 13495 19261 13504 19295
rect 13452 19252 13504 19261
rect 13728 19252 13780 19304
rect 14372 19295 14424 19304
rect 14372 19261 14381 19295
rect 14381 19261 14415 19295
rect 14415 19261 14424 19295
rect 14372 19252 14424 19261
rect 17316 19320 17368 19372
rect 20168 19456 20220 19508
rect 20996 19456 21048 19508
rect 22100 19456 22152 19508
rect 24860 19456 24912 19508
rect 19340 19320 19392 19372
rect 19984 19320 20036 19372
rect 22652 19320 22704 19372
rect 27988 19388 28040 19440
rect 25964 19363 26016 19372
rect 25964 19329 25973 19363
rect 25973 19329 26007 19363
rect 26007 19329 26016 19363
rect 25964 19320 26016 19329
rect 26148 19320 26200 19372
rect 26424 19363 26476 19372
rect 26424 19329 26433 19363
rect 26433 19329 26467 19363
rect 26467 19329 26476 19363
rect 26424 19320 26476 19329
rect 19708 19295 19760 19304
rect 19708 19261 19717 19295
rect 19717 19261 19751 19295
rect 19751 19261 19760 19295
rect 19708 19252 19760 19261
rect 20076 19252 20128 19304
rect 27344 19363 27396 19372
rect 27344 19329 27353 19363
rect 27353 19329 27387 19363
rect 27387 19329 27396 19363
rect 27344 19320 27396 19329
rect 27528 19363 27580 19372
rect 27528 19329 27536 19363
rect 27536 19329 27570 19363
rect 27570 19329 27580 19363
rect 27528 19320 27580 19329
rect 29368 19320 29420 19372
rect 28724 19252 28776 19304
rect 5908 19116 5960 19168
rect 12992 19159 13044 19168
rect 12992 19125 13001 19159
rect 13001 19125 13035 19159
rect 13035 19125 13044 19159
rect 12992 19116 13044 19125
rect 15292 19159 15344 19168
rect 15292 19125 15301 19159
rect 15301 19125 15335 19159
rect 15335 19125 15344 19159
rect 15292 19116 15344 19125
rect 19340 19116 19392 19168
rect 22836 19116 22888 19168
rect 23020 19116 23072 19168
rect 25228 19116 25280 19168
rect 25780 19159 25832 19168
rect 25780 19125 25789 19159
rect 25789 19125 25823 19159
rect 25823 19125 25832 19159
rect 25780 19116 25832 19125
rect 26608 19159 26660 19168
rect 26608 19125 26617 19159
rect 26617 19125 26651 19159
rect 26651 19125 26660 19159
rect 26608 19116 26660 19125
rect 29460 19116 29512 19168
rect 30656 19116 30708 19168
rect 4182 19014 4234 19066
rect 4246 19014 4298 19066
rect 4310 19014 4362 19066
rect 4374 19014 4426 19066
rect 4438 19014 4490 19066
rect 4502 19014 4554 19066
rect 10182 19014 10234 19066
rect 10246 19014 10298 19066
rect 10310 19014 10362 19066
rect 10374 19014 10426 19066
rect 10438 19014 10490 19066
rect 10502 19014 10554 19066
rect 16182 19014 16234 19066
rect 16246 19014 16298 19066
rect 16310 19014 16362 19066
rect 16374 19014 16426 19066
rect 16438 19014 16490 19066
rect 16502 19014 16554 19066
rect 22182 19014 22234 19066
rect 22246 19014 22298 19066
rect 22310 19014 22362 19066
rect 22374 19014 22426 19066
rect 22438 19014 22490 19066
rect 22502 19014 22554 19066
rect 28182 19014 28234 19066
rect 28246 19014 28298 19066
rect 28310 19014 28362 19066
rect 28374 19014 28426 19066
rect 28438 19014 28490 19066
rect 28502 19014 28554 19066
rect 3056 18955 3108 18964
rect 3056 18921 3065 18955
rect 3065 18921 3099 18955
rect 3099 18921 3108 18955
rect 3056 18912 3108 18921
rect 4068 18912 4120 18964
rect 5540 18912 5592 18964
rect 5908 18955 5960 18964
rect 5908 18921 5917 18955
rect 5917 18921 5951 18955
rect 5951 18921 5960 18955
rect 5908 18912 5960 18921
rect 6000 18912 6052 18964
rect 10600 18955 10652 18964
rect 10600 18921 10609 18955
rect 10609 18921 10643 18955
rect 10643 18921 10652 18955
rect 10600 18912 10652 18921
rect 4620 18776 4672 18828
rect 5172 18819 5224 18828
rect 5172 18785 5181 18819
rect 5181 18785 5215 18819
rect 5215 18785 5224 18819
rect 5172 18776 5224 18785
rect 940 18708 992 18760
rect 3148 18708 3200 18760
rect 3700 18572 3752 18624
rect 7104 18819 7156 18828
rect 7104 18785 7113 18819
rect 7113 18785 7147 18819
rect 7147 18785 7156 18819
rect 7104 18776 7156 18785
rect 7196 18776 7248 18828
rect 7748 18776 7800 18828
rect 5816 18708 5868 18760
rect 11612 18912 11664 18964
rect 11980 18912 12032 18964
rect 11520 18776 11572 18828
rect 11336 18708 11388 18760
rect 13268 18751 13320 18760
rect 13268 18717 13277 18751
rect 13277 18717 13311 18751
rect 13311 18717 13320 18751
rect 13268 18708 13320 18717
rect 14372 18912 14424 18964
rect 15384 18912 15436 18964
rect 15936 18912 15988 18964
rect 17684 18912 17736 18964
rect 16672 18844 16724 18896
rect 5540 18683 5592 18692
rect 5540 18649 5549 18683
rect 5549 18649 5583 18683
rect 5583 18649 5592 18683
rect 5540 18640 5592 18649
rect 11888 18640 11940 18692
rect 14188 18708 14240 18760
rect 14280 18708 14332 18760
rect 14464 18751 14516 18760
rect 14464 18717 14473 18751
rect 14473 18717 14507 18751
rect 14507 18717 14516 18751
rect 14464 18708 14516 18717
rect 14556 18708 14608 18760
rect 19616 18912 19668 18964
rect 20720 18912 20772 18964
rect 21180 18955 21232 18964
rect 21180 18921 21189 18955
rect 21189 18921 21223 18955
rect 21223 18921 21232 18955
rect 21180 18912 21232 18921
rect 27988 18912 28040 18964
rect 19248 18844 19300 18896
rect 22468 18844 22520 18896
rect 18236 18819 18288 18828
rect 18236 18785 18245 18819
rect 18245 18785 18279 18819
rect 18279 18785 18288 18819
rect 18236 18776 18288 18785
rect 4804 18572 4856 18624
rect 7564 18572 7616 18624
rect 13452 18572 13504 18624
rect 13912 18640 13964 18692
rect 13820 18572 13872 18624
rect 18328 18708 18380 18760
rect 21640 18819 21692 18828
rect 21640 18785 21649 18819
rect 21649 18785 21683 18819
rect 21683 18785 21692 18819
rect 21640 18776 21692 18785
rect 18052 18683 18104 18692
rect 18052 18649 18061 18683
rect 18061 18649 18095 18683
rect 18095 18649 18104 18683
rect 18052 18640 18104 18649
rect 16212 18615 16264 18624
rect 16212 18581 16221 18615
rect 16221 18581 16255 18615
rect 16255 18581 16264 18615
rect 16212 18572 16264 18581
rect 19064 18615 19116 18624
rect 19064 18581 19073 18615
rect 19073 18581 19107 18615
rect 19107 18581 19116 18615
rect 19064 18572 19116 18581
rect 21456 18708 21508 18760
rect 22100 18776 22152 18828
rect 23020 18776 23072 18828
rect 19340 18640 19392 18692
rect 19616 18572 19668 18624
rect 22744 18615 22796 18624
rect 22744 18581 22753 18615
rect 22753 18581 22787 18615
rect 22787 18581 22796 18615
rect 22744 18572 22796 18581
rect 22836 18572 22888 18624
rect 23204 18708 23256 18760
rect 26148 18708 26200 18760
rect 23020 18683 23072 18692
rect 23020 18649 23029 18683
rect 23029 18649 23063 18683
rect 23063 18649 23072 18683
rect 23020 18640 23072 18649
rect 23388 18640 23440 18692
rect 25780 18683 25832 18692
rect 25780 18649 25814 18683
rect 25814 18649 25832 18683
rect 25780 18640 25832 18649
rect 26608 18640 26660 18692
rect 27528 18708 27580 18760
rect 30564 18640 30616 18692
rect 27528 18572 27580 18624
rect 28448 18615 28500 18624
rect 28448 18581 28457 18615
rect 28457 18581 28491 18615
rect 28491 18581 28500 18615
rect 28448 18572 28500 18581
rect 4922 18470 4974 18522
rect 4986 18470 5038 18522
rect 5050 18470 5102 18522
rect 5114 18470 5166 18522
rect 5178 18470 5230 18522
rect 5242 18470 5294 18522
rect 10922 18470 10974 18522
rect 10986 18470 11038 18522
rect 11050 18470 11102 18522
rect 11114 18470 11166 18522
rect 11178 18470 11230 18522
rect 11242 18470 11294 18522
rect 16922 18470 16974 18522
rect 16986 18470 17038 18522
rect 17050 18470 17102 18522
rect 17114 18470 17166 18522
rect 17178 18470 17230 18522
rect 17242 18470 17294 18522
rect 22922 18470 22974 18522
rect 22986 18470 23038 18522
rect 23050 18470 23102 18522
rect 23114 18470 23166 18522
rect 23178 18470 23230 18522
rect 23242 18470 23294 18522
rect 28922 18470 28974 18522
rect 28986 18470 29038 18522
rect 29050 18470 29102 18522
rect 29114 18470 29166 18522
rect 29178 18470 29230 18522
rect 29242 18470 29294 18522
rect 11888 18411 11940 18420
rect 11888 18377 11897 18411
rect 11897 18377 11931 18411
rect 11931 18377 11940 18411
rect 11888 18368 11940 18377
rect 12256 18368 12308 18420
rect 12808 18368 12860 18420
rect 12900 18368 12952 18420
rect 13176 18368 13228 18420
rect 14096 18368 14148 18420
rect 14464 18368 14516 18420
rect 16212 18368 16264 18420
rect 16672 18368 16724 18420
rect 15016 18300 15068 18352
rect 18052 18368 18104 18420
rect 19064 18368 19116 18420
rect 19340 18368 19392 18420
rect 21732 18368 21784 18420
rect 25964 18411 26016 18420
rect 25964 18377 25973 18411
rect 25973 18377 26007 18411
rect 26007 18377 26016 18411
rect 25964 18368 26016 18377
rect 28448 18368 28500 18420
rect 19708 18300 19760 18352
rect 12992 18232 13044 18284
rect 8116 18164 8168 18216
rect 8484 18207 8536 18216
rect 8484 18173 8493 18207
rect 8493 18173 8527 18207
rect 8527 18173 8536 18207
rect 8484 18164 8536 18173
rect 9220 18207 9272 18216
rect 9220 18173 9229 18207
rect 9229 18173 9263 18207
rect 9263 18173 9272 18207
rect 9220 18164 9272 18173
rect 8208 18096 8260 18148
rect 12900 18164 12952 18216
rect 7288 18028 7340 18080
rect 9496 18028 9548 18080
rect 13820 18232 13872 18284
rect 14280 18275 14332 18284
rect 14280 18241 14298 18275
rect 14298 18241 14332 18275
rect 14280 18232 14332 18241
rect 14556 18207 14608 18216
rect 14556 18173 14565 18207
rect 14565 18173 14599 18207
rect 14599 18173 14608 18207
rect 14556 18164 14608 18173
rect 15660 18207 15712 18216
rect 15660 18173 15669 18207
rect 15669 18173 15703 18207
rect 15703 18173 15712 18207
rect 15660 18164 15712 18173
rect 17316 18275 17368 18284
rect 17316 18241 17325 18275
rect 17325 18241 17359 18275
rect 17359 18241 17368 18275
rect 17316 18232 17368 18241
rect 13912 18028 13964 18080
rect 14188 18028 14240 18080
rect 21180 18275 21232 18284
rect 21180 18241 21189 18275
rect 21189 18241 21223 18275
rect 21223 18241 21232 18275
rect 21180 18232 21232 18241
rect 24860 18232 24912 18284
rect 19156 18164 19208 18216
rect 20260 18207 20312 18216
rect 20260 18173 20269 18207
rect 20269 18173 20303 18207
rect 20303 18173 20312 18207
rect 20260 18164 20312 18173
rect 20352 18164 20404 18216
rect 21272 18207 21324 18216
rect 21272 18173 21281 18207
rect 21281 18173 21315 18207
rect 21315 18173 21324 18207
rect 21272 18164 21324 18173
rect 19524 18096 19576 18148
rect 18972 18028 19024 18080
rect 20076 18028 20128 18080
rect 20812 18028 20864 18080
rect 22744 18164 22796 18216
rect 28080 18300 28132 18352
rect 29368 18300 29420 18352
rect 27988 18232 28040 18284
rect 28724 18232 28776 18284
rect 21640 18096 21692 18148
rect 29736 18164 29788 18216
rect 29552 18096 29604 18148
rect 26424 18028 26476 18080
rect 29460 18028 29512 18080
rect 4182 17926 4234 17978
rect 4246 17926 4298 17978
rect 4310 17926 4362 17978
rect 4374 17926 4426 17978
rect 4438 17926 4490 17978
rect 4502 17926 4554 17978
rect 10182 17926 10234 17978
rect 10246 17926 10298 17978
rect 10310 17926 10362 17978
rect 10374 17926 10426 17978
rect 10438 17926 10490 17978
rect 10502 17926 10554 17978
rect 16182 17926 16234 17978
rect 16246 17926 16298 17978
rect 16310 17926 16362 17978
rect 16374 17926 16426 17978
rect 16438 17926 16490 17978
rect 16502 17926 16554 17978
rect 22182 17926 22234 17978
rect 22246 17926 22298 17978
rect 22310 17926 22362 17978
rect 22374 17926 22426 17978
rect 22438 17926 22490 17978
rect 22502 17926 22554 17978
rect 28182 17926 28234 17978
rect 28246 17926 28298 17978
rect 28310 17926 28362 17978
rect 28374 17926 28426 17978
rect 28438 17926 28490 17978
rect 28502 17926 28554 17978
rect 8852 17824 8904 17876
rect 9220 17824 9272 17876
rect 13268 17824 13320 17876
rect 14280 17867 14332 17876
rect 14280 17833 14289 17867
rect 14289 17833 14323 17867
rect 14323 17833 14332 17867
rect 14280 17824 14332 17833
rect 15384 17824 15436 17876
rect 5816 17756 5868 17808
rect 15292 17756 15344 17808
rect 21180 17824 21232 17876
rect 21272 17824 21324 17876
rect 30196 17756 30248 17808
rect 12624 17688 12676 17740
rect 6920 17620 6972 17672
rect 7288 17663 7340 17672
rect 7288 17629 7322 17663
rect 7322 17629 7340 17663
rect 7288 17620 7340 17629
rect 12164 17663 12216 17672
rect 12164 17629 12173 17663
rect 12173 17629 12207 17663
rect 12207 17629 12216 17663
rect 12164 17620 12216 17629
rect 12440 17663 12492 17672
rect 12440 17629 12449 17663
rect 12449 17629 12483 17663
rect 12483 17629 12492 17663
rect 12440 17620 12492 17629
rect 12532 17663 12584 17672
rect 12532 17629 12541 17663
rect 12541 17629 12575 17663
rect 12575 17629 12584 17663
rect 12532 17620 12584 17629
rect 5724 17552 5776 17604
rect 6092 17595 6144 17604
rect 6092 17561 6101 17595
rect 6101 17561 6135 17595
rect 6135 17561 6144 17595
rect 6092 17552 6144 17561
rect 12348 17595 12400 17604
rect 12348 17561 12357 17595
rect 12357 17561 12391 17595
rect 12391 17561 12400 17595
rect 12348 17552 12400 17561
rect 4804 17484 4856 17536
rect 5356 17484 5408 17536
rect 6368 17527 6420 17536
rect 6368 17493 6377 17527
rect 6377 17493 6411 17527
rect 6411 17493 6420 17527
rect 6368 17484 6420 17493
rect 13544 17527 13596 17536
rect 13544 17493 13553 17527
rect 13553 17493 13587 17527
rect 13587 17493 13596 17527
rect 13544 17484 13596 17493
rect 14004 17484 14056 17536
rect 14924 17688 14976 17740
rect 15476 17688 15528 17740
rect 16488 17663 16540 17672
rect 16488 17629 16497 17663
rect 16497 17629 16531 17663
rect 16531 17629 16540 17663
rect 16488 17620 16540 17629
rect 18420 17595 18472 17604
rect 18420 17561 18429 17595
rect 18429 17561 18463 17595
rect 18463 17561 18472 17595
rect 18420 17552 18472 17561
rect 19340 17620 19392 17672
rect 19984 17688 20036 17740
rect 26884 17688 26936 17740
rect 29368 17731 29420 17740
rect 29368 17697 29377 17731
rect 29377 17697 29411 17731
rect 29411 17697 29420 17731
rect 29368 17688 29420 17697
rect 29736 17731 29788 17740
rect 29736 17697 29745 17731
rect 29745 17697 29779 17731
rect 29779 17697 29788 17731
rect 29736 17688 29788 17697
rect 19524 17663 19576 17672
rect 19524 17629 19533 17663
rect 19533 17629 19567 17663
rect 19567 17629 19576 17663
rect 19524 17620 19576 17629
rect 19800 17620 19852 17672
rect 20444 17663 20496 17672
rect 20444 17629 20453 17663
rect 20453 17629 20487 17663
rect 20487 17629 20496 17663
rect 20444 17620 20496 17629
rect 20720 17663 20772 17672
rect 20720 17629 20729 17663
rect 20729 17629 20763 17663
rect 20763 17629 20772 17663
rect 20720 17620 20772 17629
rect 20904 17620 20956 17672
rect 21548 17620 21600 17672
rect 23940 17620 23992 17672
rect 20352 17552 20404 17604
rect 21732 17552 21784 17604
rect 15016 17484 15068 17536
rect 15844 17484 15896 17536
rect 17868 17484 17920 17536
rect 19340 17484 19392 17536
rect 25044 17527 25096 17536
rect 25044 17493 25053 17527
rect 25053 17493 25087 17527
rect 25087 17493 25096 17527
rect 25044 17484 25096 17493
rect 28724 17527 28776 17536
rect 28724 17493 28733 17527
rect 28733 17493 28767 17527
rect 28767 17493 28776 17527
rect 28724 17484 28776 17493
rect 28816 17484 28868 17536
rect 29920 17527 29972 17536
rect 29920 17493 29929 17527
rect 29929 17493 29963 17527
rect 29963 17493 29972 17527
rect 29920 17484 29972 17493
rect 4922 17382 4974 17434
rect 4986 17382 5038 17434
rect 5050 17382 5102 17434
rect 5114 17382 5166 17434
rect 5178 17382 5230 17434
rect 5242 17382 5294 17434
rect 10922 17382 10974 17434
rect 10986 17382 11038 17434
rect 11050 17382 11102 17434
rect 11114 17382 11166 17434
rect 11178 17382 11230 17434
rect 11242 17382 11294 17434
rect 16922 17382 16974 17434
rect 16986 17382 17038 17434
rect 17050 17382 17102 17434
rect 17114 17382 17166 17434
rect 17178 17382 17230 17434
rect 17242 17382 17294 17434
rect 22922 17382 22974 17434
rect 22986 17382 23038 17434
rect 23050 17382 23102 17434
rect 23114 17382 23166 17434
rect 23178 17382 23230 17434
rect 23242 17382 23294 17434
rect 28922 17382 28974 17434
rect 28986 17382 29038 17434
rect 29050 17382 29102 17434
rect 29114 17382 29166 17434
rect 29178 17382 29230 17434
rect 29242 17382 29294 17434
rect 4804 17323 4856 17332
rect 4804 17289 4813 17323
rect 4813 17289 4847 17323
rect 4847 17289 4856 17323
rect 4804 17280 4856 17289
rect 5356 17280 5408 17332
rect 6368 17280 6420 17332
rect 7012 17212 7064 17264
rect 8852 17255 8904 17264
rect 8852 17221 8861 17255
rect 8861 17221 8895 17255
rect 8895 17221 8904 17255
rect 8852 17212 8904 17221
rect 3516 17144 3568 17196
rect 3976 17144 4028 17196
rect 8760 17187 8812 17196
rect 8760 17153 8769 17187
rect 8769 17153 8803 17187
rect 8803 17153 8812 17187
rect 8760 17144 8812 17153
rect 13544 17280 13596 17332
rect 15844 17280 15896 17332
rect 15200 17212 15252 17264
rect 15752 17212 15804 17264
rect 16488 17280 16540 17332
rect 19340 17280 19392 17332
rect 25044 17280 25096 17332
rect 26240 17280 26292 17332
rect 27160 17280 27212 17332
rect 28724 17280 28776 17332
rect 28816 17280 28868 17332
rect 29184 17280 29236 17332
rect 29368 17280 29420 17332
rect 29920 17280 29972 17332
rect 19800 17212 19852 17264
rect 20352 17212 20404 17264
rect 10600 17144 10652 17196
rect 14004 17144 14056 17196
rect 14188 17144 14240 17196
rect 17316 17144 17368 17196
rect 18236 17144 18288 17196
rect 22652 17144 22704 17196
rect 4620 17076 4672 17128
rect 5356 17119 5408 17128
rect 5356 17085 5365 17119
rect 5365 17085 5399 17119
rect 5399 17085 5408 17119
rect 5356 17076 5408 17085
rect 4896 16983 4948 16992
rect 4896 16949 4905 16983
rect 4905 16949 4939 16983
rect 4939 16949 4948 16983
rect 4896 16940 4948 16949
rect 13912 17119 13964 17128
rect 13912 17085 13921 17119
rect 13921 17085 13955 17119
rect 13955 17085 13964 17119
rect 13912 17076 13964 17085
rect 23572 17119 23624 17128
rect 23572 17085 23581 17119
rect 23581 17085 23615 17119
rect 23615 17085 23624 17119
rect 23572 17076 23624 17085
rect 23848 17187 23900 17196
rect 23848 17153 23857 17187
rect 23857 17153 23891 17187
rect 23891 17153 23900 17187
rect 23848 17144 23900 17153
rect 23940 17144 23992 17196
rect 26056 17144 26108 17196
rect 26240 17187 26292 17196
rect 26240 17153 26249 17187
rect 26249 17153 26283 17187
rect 26283 17153 26292 17187
rect 26240 17144 26292 17153
rect 26884 17212 26936 17264
rect 27620 17212 27672 17264
rect 29092 17212 29144 17264
rect 29460 17212 29512 17264
rect 9128 17008 9180 17060
rect 19892 17008 19944 17060
rect 20260 17008 20312 17060
rect 25688 17008 25740 17060
rect 25872 17119 25924 17128
rect 25872 17085 25881 17119
rect 25881 17085 25915 17119
rect 25915 17085 25924 17119
rect 29828 17212 29880 17264
rect 28080 17144 28132 17196
rect 29644 17144 29696 17196
rect 30564 17144 30616 17196
rect 25872 17076 25924 17085
rect 26240 17008 26292 17060
rect 6920 16940 6972 16992
rect 7840 16940 7892 16992
rect 8024 16983 8076 16992
rect 8024 16949 8033 16983
rect 8033 16949 8067 16983
rect 8067 16949 8076 16983
rect 8024 16940 8076 16949
rect 9036 16940 9088 16992
rect 9680 16940 9732 16992
rect 10048 16940 10100 16992
rect 12072 16940 12124 16992
rect 22100 16940 22152 16992
rect 22744 16940 22796 16992
rect 24032 16983 24084 16992
rect 24032 16949 24041 16983
rect 24041 16949 24075 16983
rect 24075 16949 24084 16983
rect 24032 16940 24084 16949
rect 25320 16983 25372 16992
rect 25320 16949 25329 16983
rect 25329 16949 25363 16983
rect 25363 16949 25372 16983
rect 25320 16940 25372 16949
rect 25780 16940 25832 16992
rect 30932 17119 30984 17128
rect 30932 17085 30941 17119
rect 30941 17085 30975 17119
rect 30975 17085 30984 17119
rect 30932 17076 30984 17085
rect 4182 16838 4234 16890
rect 4246 16838 4298 16890
rect 4310 16838 4362 16890
rect 4374 16838 4426 16890
rect 4438 16838 4490 16890
rect 4502 16838 4554 16890
rect 10182 16838 10234 16890
rect 10246 16838 10298 16890
rect 10310 16838 10362 16890
rect 10374 16838 10426 16890
rect 10438 16838 10490 16890
rect 10502 16838 10554 16890
rect 16182 16838 16234 16890
rect 16246 16838 16298 16890
rect 16310 16838 16362 16890
rect 16374 16838 16426 16890
rect 16438 16838 16490 16890
rect 16502 16838 16554 16890
rect 22182 16838 22234 16890
rect 22246 16838 22298 16890
rect 22310 16838 22362 16890
rect 22374 16838 22426 16890
rect 22438 16838 22490 16890
rect 22502 16838 22554 16890
rect 28182 16838 28234 16890
rect 28246 16838 28298 16890
rect 28310 16838 28362 16890
rect 28374 16838 28426 16890
rect 28438 16838 28490 16890
rect 28502 16838 28554 16890
rect 3516 16736 3568 16788
rect 3976 16736 4028 16788
rect 7012 16736 7064 16788
rect 8760 16736 8812 16788
rect 5356 16668 5408 16720
rect 3424 16575 3476 16584
rect 3424 16541 3433 16575
rect 3433 16541 3467 16575
rect 3467 16541 3476 16575
rect 3424 16532 3476 16541
rect 4896 16532 4948 16584
rect 4620 16464 4672 16516
rect 6092 16600 6144 16652
rect 9128 16668 9180 16720
rect 11704 16668 11756 16720
rect 12072 16736 12124 16788
rect 13084 16736 13136 16788
rect 15200 16736 15252 16788
rect 18236 16779 18288 16788
rect 18236 16745 18245 16779
rect 18245 16745 18279 16779
rect 18279 16745 18288 16779
rect 18236 16736 18288 16745
rect 19156 16736 19208 16788
rect 6828 16532 6880 16584
rect 7380 16600 7432 16652
rect 7840 16600 7892 16652
rect 14648 16668 14700 16720
rect 14188 16600 14240 16652
rect 14372 16600 14424 16652
rect 23848 16736 23900 16788
rect 25872 16736 25924 16788
rect 28632 16736 28684 16788
rect 27160 16668 27212 16720
rect 29460 16736 29512 16788
rect 29920 16736 29972 16788
rect 8024 16532 8076 16584
rect 10048 16575 10100 16584
rect 10048 16541 10082 16575
rect 10082 16541 10100 16575
rect 10048 16532 10100 16541
rect 18972 16532 19024 16584
rect 21548 16532 21600 16584
rect 22100 16575 22152 16584
rect 22100 16541 22134 16575
rect 22134 16541 22152 16575
rect 22100 16532 22152 16541
rect 23848 16532 23900 16584
rect 24032 16532 24084 16584
rect 29092 16600 29144 16652
rect 29184 16600 29236 16652
rect 25596 16532 25648 16584
rect 25688 16532 25740 16584
rect 28908 16575 28960 16584
rect 28908 16541 28912 16575
rect 28912 16541 28946 16575
rect 28946 16541 28960 16575
rect 28908 16532 28960 16541
rect 29460 16532 29512 16584
rect 30196 16532 30248 16584
rect 30932 16532 30984 16584
rect 25320 16464 25372 16516
rect 30656 16464 30708 16516
rect 9588 16396 9640 16448
rect 11336 16396 11388 16448
rect 23388 16396 23440 16448
rect 25872 16439 25924 16448
rect 25872 16405 25881 16439
rect 25881 16405 25915 16439
rect 25915 16405 25924 16439
rect 25872 16396 25924 16405
rect 4922 16294 4974 16346
rect 4986 16294 5038 16346
rect 5050 16294 5102 16346
rect 5114 16294 5166 16346
rect 5178 16294 5230 16346
rect 5242 16294 5294 16346
rect 10922 16294 10974 16346
rect 10986 16294 11038 16346
rect 11050 16294 11102 16346
rect 11114 16294 11166 16346
rect 11178 16294 11230 16346
rect 11242 16294 11294 16346
rect 16922 16294 16974 16346
rect 16986 16294 17038 16346
rect 17050 16294 17102 16346
rect 17114 16294 17166 16346
rect 17178 16294 17230 16346
rect 17242 16294 17294 16346
rect 22922 16294 22974 16346
rect 22986 16294 23038 16346
rect 23050 16294 23102 16346
rect 23114 16294 23166 16346
rect 23178 16294 23230 16346
rect 23242 16294 23294 16346
rect 28922 16294 28974 16346
rect 28986 16294 29038 16346
rect 29050 16294 29102 16346
rect 29114 16294 29166 16346
rect 29178 16294 29230 16346
rect 29242 16294 29294 16346
rect 3424 16192 3476 16244
rect 4620 16235 4672 16244
rect 4620 16201 4629 16235
rect 4629 16201 4663 16235
rect 4663 16201 4672 16235
rect 4620 16192 4672 16201
rect 5356 16192 5408 16244
rect 9496 16192 9548 16244
rect 10600 16192 10652 16244
rect 11336 16192 11388 16244
rect 8944 16099 8996 16108
rect 8944 16065 8953 16099
rect 8953 16065 8987 16099
rect 8987 16065 8996 16099
rect 8944 16056 8996 16065
rect 9036 16099 9088 16108
rect 9036 16065 9046 16099
rect 9046 16065 9080 16099
rect 9080 16065 9088 16099
rect 9036 16056 9088 16065
rect 9312 16099 9364 16108
rect 9312 16065 9321 16099
rect 9321 16065 9355 16099
rect 9355 16065 9364 16099
rect 9312 16056 9364 16065
rect 9588 16056 9640 16108
rect 9680 16056 9732 16108
rect 11704 16167 11756 16176
rect 11704 16133 11713 16167
rect 11713 16133 11747 16167
rect 11747 16133 11756 16167
rect 11704 16124 11756 16133
rect 11796 16056 11848 16108
rect 15200 16099 15252 16108
rect 15200 16065 15209 16099
rect 15209 16065 15243 16099
rect 15243 16065 15252 16099
rect 15200 16056 15252 16065
rect 15752 16056 15804 16108
rect 21732 16192 21784 16244
rect 4804 16031 4856 16040
rect 4804 15997 4813 16031
rect 4813 15997 4847 16031
rect 4847 15997 4856 16031
rect 4804 15988 4856 15997
rect 10692 15988 10744 16040
rect 10600 15852 10652 15904
rect 10784 15920 10836 15972
rect 21364 15988 21416 16040
rect 15568 15852 15620 15904
rect 17960 15852 18012 15904
rect 21180 15852 21232 15904
rect 21548 15988 21600 16040
rect 22100 15852 22152 15904
rect 23204 16056 23256 16108
rect 23388 16124 23440 16176
rect 23572 16167 23624 16176
rect 23572 16133 23581 16167
rect 23581 16133 23615 16167
rect 23615 16133 23624 16167
rect 23572 16124 23624 16133
rect 25872 16124 25924 16176
rect 26056 16192 26108 16244
rect 27620 16192 27672 16244
rect 25596 15988 25648 16040
rect 25780 16099 25832 16108
rect 25780 16065 25789 16099
rect 25789 16065 25823 16099
rect 25823 16065 25832 16099
rect 25780 16056 25832 16065
rect 26148 16056 26200 16108
rect 27160 16056 27212 16108
rect 27068 16031 27120 16040
rect 27068 15997 27077 16031
rect 27077 15997 27111 16031
rect 27111 15997 27120 16031
rect 27068 15988 27120 15997
rect 27896 15988 27948 16040
rect 23572 15920 23624 15972
rect 23940 15895 23992 15904
rect 23940 15861 23949 15895
rect 23949 15861 23983 15895
rect 23983 15861 23992 15895
rect 23940 15852 23992 15861
rect 26240 15852 26292 15904
rect 26516 15895 26568 15904
rect 26516 15861 26525 15895
rect 26525 15861 26559 15895
rect 26559 15861 26568 15895
rect 26516 15852 26568 15861
rect 27712 15895 27764 15904
rect 27712 15861 27721 15895
rect 27721 15861 27755 15895
rect 27755 15861 27764 15895
rect 27712 15852 27764 15861
rect 4182 15750 4234 15802
rect 4246 15750 4298 15802
rect 4310 15750 4362 15802
rect 4374 15750 4426 15802
rect 4438 15750 4490 15802
rect 4502 15750 4554 15802
rect 10182 15750 10234 15802
rect 10246 15750 10298 15802
rect 10310 15750 10362 15802
rect 10374 15750 10426 15802
rect 10438 15750 10490 15802
rect 10502 15750 10554 15802
rect 16182 15750 16234 15802
rect 16246 15750 16298 15802
rect 16310 15750 16362 15802
rect 16374 15750 16426 15802
rect 16438 15750 16490 15802
rect 16502 15750 16554 15802
rect 22182 15750 22234 15802
rect 22246 15750 22298 15802
rect 22310 15750 22362 15802
rect 22374 15750 22426 15802
rect 22438 15750 22490 15802
rect 22502 15750 22554 15802
rect 28182 15750 28234 15802
rect 28246 15750 28298 15802
rect 28310 15750 28362 15802
rect 28374 15750 28426 15802
rect 28438 15750 28490 15802
rect 28502 15750 28554 15802
rect 8944 15648 8996 15700
rect 9312 15648 9364 15700
rect 8760 15623 8812 15632
rect 8760 15589 8769 15623
rect 8769 15589 8803 15623
rect 8803 15589 8812 15623
rect 8760 15580 8812 15589
rect 15568 15648 15620 15700
rect 22376 15648 22428 15700
rect 22652 15648 22704 15700
rect 23388 15648 23440 15700
rect 26148 15691 26200 15700
rect 26148 15657 26157 15691
rect 26157 15657 26191 15691
rect 26191 15657 26200 15691
rect 26148 15648 26200 15657
rect 27712 15648 27764 15700
rect 7196 15487 7248 15496
rect 7196 15453 7205 15487
rect 7205 15453 7239 15487
rect 7239 15453 7248 15487
rect 7196 15444 7248 15453
rect 7840 15444 7892 15496
rect 8300 15444 8352 15496
rect 8576 15487 8628 15496
rect 8576 15453 8585 15487
rect 8585 15453 8619 15487
rect 8619 15453 8628 15487
rect 8576 15444 8628 15453
rect 6644 15351 6696 15360
rect 6644 15317 6653 15351
rect 6653 15317 6687 15351
rect 6687 15317 6696 15351
rect 6644 15308 6696 15317
rect 8760 15376 8812 15428
rect 10416 15487 10468 15496
rect 10416 15453 10425 15487
rect 10425 15453 10459 15487
rect 10459 15453 10468 15487
rect 10416 15444 10468 15453
rect 11980 15487 12032 15496
rect 11980 15453 11989 15487
rect 11989 15453 12023 15487
rect 12023 15453 12032 15487
rect 11980 15444 12032 15453
rect 12808 15444 12860 15496
rect 17776 15487 17828 15496
rect 17776 15453 17785 15487
rect 17785 15453 17819 15487
rect 17819 15453 17828 15487
rect 17776 15444 17828 15453
rect 18144 15487 18196 15496
rect 18144 15453 18153 15487
rect 18153 15453 18187 15487
rect 18187 15453 18196 15487
rect 18144 15444 18196 15453
rect 18236 15444 18288 15496
rect 20076 15444 20128 15496
rect 21732 15580 21784 15632
rect 22560 15580 22612 15632
rect 23204 15580 23256 15632
rect 12532 15376 12584 15428
rect 18052 15376 18104 15428
rect 19708 15376 19760 15428
rect 20904 15444 20956 15496
rect 20996 15444 21048 15496
rect 22928 15555 22980 15564
rect 22928 15521 22937 15555
rect 22937 15521 22971 15555
rect 22971 15521 22980 15555
rect 22928 15512 22980 15521
rect 23020 15555 23072 15564
rect 23020 15521 23029 15555
rect 23029 15521 23063 15555
rect 23063 15521 23072 15555
rect 23020 15512 23072 15521
rect 25228 15512 25280 15564
rect 22468 15444 22520 15496
rect 25596 15444 25648 15496
rect 27528 15444 27580 15496
rect 23940 15376 23992 15428
rect 26056 15376 26108 15428
rect 26516 15419 26568 15428
rect 26516 15385 26550 15419
rect 26550 15385 26568 15419
rect 26516 15376 26568 15385
rect 12348 15308 12400 15360
rect 12900 15308 12952 15360
rect 17592 15351 17644 15360
rect 17592 15317 17601 15351
rect 17601 15317 17635 15351
rect 17635 15317 17644 15351
rect 17592 15308 17644 15317
rect 18512 15308 18564 15360
rect 18604 15351 18656 15360
rect 18604 15317 18613 15351
rect 18613 15317 18647 15351
rect 18647 15317 18656 15351
rect 18604 15308 18656 15317
rect 20904 15308 20956 15360
rect 21180 15308 21232 15360
rect 23020 15308 23072 15360
rect 27620 15351 27672 15360
rect 27620 15317 27629 15351
rect 27629 15317 27663 15351
rect 27663 15317 27672 15351
rect 27620 15308 27672 15317
rect 28264 15308 28316 15360
rect 4922 15206 4974 15258
rect 4986 15206 5038 15258
rect 5050 15206 5102 15258
rect 5114 15206 5166 15258
rect 5178 15206 5230 15258
rect 5242 15206 5294 15258
rect 10922 15206 10974 15258
rect 10986 15206 11038 15258
rect 11050 15206 11102 15258
rect 11114 15206 11166 15258
rect 11178 15206 11230 15258
rect 11242 15206 11294 15258
rect 16922 15206 16974 15258
rect 16986 15206 17038 15258
rect 17050 15206 17102 15258
rect 17114 15206 17166 15258
rect 17178 15206 17230 15258
rect 17242 15206 17294 15258
rect 22922 15206 22974 15258
rect 22986 15206 23038 15258
rect 23050 15206 23102 15258
rect 23114 15206 23166 15258
rect 23178 15206 23230 15258
rect 23242 15206 23294 15258
rect 28922 15206 28974 15258
rect 28986 15206 29038 15258
rect 29050 15206 29102 15258
rect 29114 15206 29166 15258
rect 29178 15206 29230 15258
rect 29242 15206 29294 15258
rect 6644 15104 6696 15156
rect 6828 15147 6880 15156
rect 6828 15113 6837 15147
rect 6837 15113 6871 15147
rect 6871 15113 6880 15147
rect 6828 15104 6880 15113
rect 8116 15104 8168 15156
rect 8576 15104 8628 15156
rect 10416 15104 10468 15156
rect 12624 15104 12676 15156
rect 18972 15104 19024 15156
rect 10692 15036 10744 15088
rect 12440 15079 12492 15088
rect 12440 15045 12474 15079
rect 12474 15045 12492 15079
rect 12440 15036 12492 15045
rect 1676 14900 1728 14952
rect 4068 14900 4120 14952
rect 7932 15011 7984 15020
rect 7932 14977 7941 15011
rect 7941 14977 7975 15011
rect 7975 14977 7984 15011
rect 7932 14968 7984 14977
rect 14648 15036 14700 15088
rect 4804 14900 4856 14952
rect 7104 14900 7156 14952
rect 8208 14943 8260 14952
rect 8208 14909 8217 14943
rect 8217 14909 8251 14943
rect 8251 14909 8260 14943
rect 8208 14900 8260 14909
rect 13268 14968 13320 15020
rect 18328 15036 18380 15088
rect 17592 15011 17644 15020
rect 17592 14977 17626 15011
rect 17626 14977 17644 15011
rect 17592 14968 17644 14977
rect 18512 14968 18564 15020
rect 21548 15036 21600 15088
rect 22100 15104 22152 15156
rect 22744 15104 22796 15156
rect 26240 15147 26292 15156
rect 26240 15113 26249 15147
rect 26249 15113 26283 15147
rect 26283 15113 26292 15147
rect 26240 15104 26292 15113
rect 2688 14807 2740 14816
rect 2688 14773 2697 14807
rect 2697 14773 2731 14807
rect 2731 14773 2740 14807
rect 2688 14764 2740 14773
rect 3516 14764 3568 14816
rect 4620 14764 4672 14816
rect 6368 14807 6420 14816
rect 6368 14773 6377 14807
rect 6377 14773 6411 14807
rect 6411 14773 6420 14807
rect 6368 14764 6420 14773
rect 7564 14807 7616 14816
rect 7564 14773 7573 14807
rect 7573 14773 7607 14807
rect 7607 14773 7616 14807
rect 7564 14764 7616 14773
rect 12532 14764 12584 14816
rect 13452 14764 13504 14816
rect 21272 14968 21324 15020
rect 22376 14968 22428 15020
rect 23940 14968 23992 15020
rect 20996 14943 21048 14952
rect 20996 14909 21005 14943
rect 21005 14909 21039 14943
rect 21039 14909 21048 14943
rect 20996 14900 21048 14909
rect 20168 14875 20220 14884
rect 20168 14841 20177 14875
rect 20177 14841 20211 14875
rect 20211 14841 20220 14875
rect 20168 14832 20220 14841
rect 21364 14832 21416 14884
rect 13636 14807 13688 14816
rect 13636 14773 13645 14807
rect 13645 14773 13679 14807
rect 13679 14773 13688 14807
rect 13636 14764 13688 14773
rect 14372 14807 14424 14816
rect 14372 14773 14381 14807
rect 14381 14773 14415 14807
rect 14415 14773 14424 14807
rect 14372 14764 14424 14773
rect 20076 14764 20128 14816
rect 20260 14807 20312 14816
rect 20260 14773 20269 14807
rect 20269 14773 20303 14807
rect 20303 14773 20312 14807
rect 20260 14764 20312 14773
rect 20812 14764 20864 14816
rect 21640 14807 21692 14816
rect 21640 14773 21649 14807
rect 21649 14773 21683 14807
rect 21683 14773 21692 14807
rect 21640 14764 21692 14773
rect 27896 15104 27948 15156
rect 27528 15036 27580 15088
rect 26424 15011 26476 15020
rect 26424 14977 26433 15011
rect 26433 14977 26467 15011
rect 26467 14977 26476 15011
rect 26424 14968 26476 14977
rect 26700 14968 26752 15020
rect 27620 14968 27672 15020
rect 28264 14968 28316 15020
rect 28632 14968 28684 15020
rect 31208 14764 31260 14816
rect 4182 14662 4234 14714
rect 4246 14662 4298 14714
rect 4310 14662 4362 14714
rect 4374 14662 4426 14714
rect 4438 14662 4490 14714
rect 4502 14662 4554 14714
rect 10182 14662 10234 14714
rect 10246 14662 10298 14714
rect 10310 14662 10362 14714
rect 10374 14662 10426 14714
rect 10438 14662 10490 14714
rect 10502 14662 10554 14714
rect 16182 14662 16234 14714
rect 16246 14662 16298 14714
rect 16310 14662 16362 14714
rect 16374 14662 16426 14714
rect 16438 14662 16490 14714
rect 16502 14662 16554 14714
rect 22182 14662 22234 14714
rect 22246 14662 22298 14714
rect 22310 14662 22362 14714
rect 22374 14662 22426 14714
rect 22438 14662 22490 14714
rect 22502 14662 22554 14714
rect 28182 14662 28234 14714
rect 28246 14662 28298 14714
rect 28310 14662 28362 14714
rect 28374 14662 28426 14714
rect 28438 14662 28490 14714
rect 28502 14662 28554 14714
rect 7196 14560 7248 14612
rect 7840 14603 7892 14612
rect 7840 14569 7849 14603
rect 7849 14569 7883 14603
rect 7883 14569 7892 14603
rect 7840 14560 7892 14569
rect 7932 14603 7984 14612
rect 7932 14569 7941 14603
rect 7941 14569 7975 14603
rect 7975 14569 7984 14603
rect 7932 14560 7984 14569
rect 12440 14603 12492 14612
rect 12440 14569 12449 14603
rect 12449 14569 12483 14603
rect 12483 14569 12492 14603
rect 12440 14560 12492 14569
rect 13636 14560 13688 14612
rect 17776 14560 17828 14612
rect 17960 14560 18012 14612
rect 18144 14560 18196 14612
rect 4712 14424 4764 14476
rect 8300 14356 8352 14408
rect 3240 14288 3292 14340
rect 3516 14288 3568 14340
rect 2320 14220 2372 14272
rect 3608 14263 3660 14272
rect 3608 14229 3617 14263
rect 3617 14229 3651 14263
rect 3651 14229 3660 14263
rect 3608 14220 3660 14229
rect 3792 14263 3844 14272
rect 3792 14229 3801 14263
rect 3801 14229 3835 14263
rect 3835 14229 3844 14263
rect 3792 14220 3844 14229
rect 4160 14263 4212 14272
rect 4160 14229 4169 14263
rect 4169 14229 4203 14263
rect 4203 14229 4212 14263
rect 4160 14220 4212 14229
rect 6000 14288 6052 14340
rect 7012 14288 7064 14340
rect 7840 14288 7892 14340
rect 13360 14467 13412 14476
rect 13360 14433 13369 14467
rect 13369 14433 13403 14467
rect 13403 14433 13412 14467
rect 13360 14424 13412 14433
rect 13544 14424 13596 14476
rect 16028 14535 16080 14544
rect 16028 14501 16037 14535
rect 16037 14501 16071 14535
rect 16071 14501 16080 14535
rect 16028 14492 16080 14501
rect 13728 14399 13780 14408
rect 13728 14365 13737 14399
rect 13737 14365 13771 14399
rect 13771 14365 13780 14399
rect 13728 14356 13780 14365
rect 14096 14356 14148 14408
rect 14740 14356 14792 14408
rect 10784 14220 10836 14272
rect 14464 14288 14516 14340
rect 11888 14220 11940 14272
rect 12808 14220 12860 14272
rect 13544 14263 13596 14272
rect 13544 14229 13553 14263
rect 13553 14229 13587 14263
rect 13587 14229 13596 14263
rect 13544 14220 13596 14229
rect 16120 14263 16172 14272
rect 16120 14229 16129 14263
rect 16129 14229 16163 14263
rect 16163 14229 16172 14263
rect 16120 14220 16172 14229
rect 16672 14220 16724 14272
rect 18512 14467 18564 14476
rect 18512 14433 18521 14467
rect 18521 14433 18555 14467
rect 18555 14433 18564 14467
rect 18512 14424 18564 14433
rect 19156 14424 19208 14476
rect 18144 14356 18196 14408
rect 18236 14356 18288 14408
rect 20260 14560 20312 14612
rect 20904 14560 20956 14612
rect 21732 14560 21784 14612
rect 19892 14467 19944 14476
rect 19892 14433 19901 14467
rect 19901 14433 19935 14467
rect 19935 14433 19944 14467
rect 19892 14424 19944 14433
rect 21364 14399 21416 14408
rect 21364 14365 21382 14399
rect 21382 14365 21416 14399
rect 21364 14356 21416 14365
rect 21548 14356 21600 14408
rect 18052 14220 18104 14272
rect 20996 14220 21048 14272
rect 21088 14220 21140 14272
rect 4922 14118 4974 14170
rect 4986 14118 5038 14170
rect 5050 14118 5102 14170
rect 5114 14118 5166 14170
rect 5178 14118 5230 14170
rect 5242 14118 5294 14170
rect 10922 14118 10974 14170
rect 10986 14118 11038 14170
rect 11050 14118 11102 14170
rect 11114 14118 11166 14170
rect 11178 14118 11230 14170
rect 11242 14118 11294 14170
rect 16922 14118 16974 14170
rect 16986 14118 17038 14170
rect 17050 14118 17102 14170
rect 17114 14118 17166 14170
rect 17178 14118 17230 14170
rect 17242 14118 17294 14170
rect 22922 14118 22974 14170
rect 22986 14118 23038 14170
rect 23050 14118 23102 14170
rect 23114 14118 23166 14170
rect 23178 14118 23230 14170
rect 23242 14118 23294 14170
rect 28922 14118 28974 14170
rect 28986 14118 29038 14170
rect 29050 14118 29102 14170
rect 29114 14118 29166 14170
rect 29178 14118 29230 14170
rect 29242 14118 29294 14170
rect 2688 14016 2740 14068
rect 3608 14016 3660 14068
rect 2320 13923 2372 13932
rect 2320 13889 2329 13923
rect 2329 13889 2363 13923
rect 2363 13889 2372 13923
rect 2320 13880 2372 13889
rect 4160 14016 4212 14068
rect 4620 13948 4672 14000
rect 5356 14016 5408 14068
rect 5816 14016 5868 14068
rect 6000 14059 6052 14068
rect 6000 14025 6009 14059
rect 6009 14025 6043 14059
rect 6043 14025 6052 14059
rect 6000 14016 6052 14025
rect 6368 14016 6420 14068
rect 7012 14059 7064 14068
rect 7012 14025 7021 14059
rect 7021 14025 7055 14059
rect 7055 14025 7064 14059
rect 7012 14016 7064 14025
rect 7564 14016 7616 14068
rect 10784 14016 10836 14068
rect 5448 13948 5500 14000
rect 5724 13948 5776 14000
rect 11980 14016 12032 14068
rect 13084 14016 13136 14068
rect 13268 14016 13320 14068
rect 13728 14016 13780 14068
rect 14372 14016 14424 14068
rect 14464 14016 14516 14068
rect 14740 14016 14792 14068
rect 16120 14016 16172 14068
rect 18328 14016 18380 14068
rect 19708 14059 19760 14068
rect 19708 14025 19717 14059
rect 19717 14025 19751 14059
rect 19751 14025 19760 14059
rect 19708 14016 19760 14025
rect 13544 13991 13596 14000
rect 13544 13957 13562 13991
rect 13562 13957 13596 13991
rect 13544 13948 13596 13957
rect 11888 13812 11940 13864
rect 12072 13855 12124 13864
rect 12072 13821 12081 13855
rect 12081 13821 12115 13855
rect 12115 13821 12124 13855
rect 12072 13812 12124 13821
rect 14096 13812 14148 13864
rect 14464 13855 14516 13864
rect 14464 13821 14473 13855
rect 14473 13821 14507 13855
rect 14507 13821 14516 13855
rect 14464 13812 14516 13821
rect 15384 13855 15436 13864
rect 15384 13821 15393 13855
rect 15393 13821 15427 13855
rect 15427 13821 15436 13855
rect 15384 13812 15436 13821
rect 15752 13923 15804 13932
rect 15752 13889 15761 13923
rect 15761 13889 15795 13923
rect 15795 13889 15804 13923
rect 15752 13880 15804 13889
rect 16028 13948 16080 14000
rect 16672 13923 16724 13932
rect 16672 13889 16681 13923
rect 16681 13889 16715 13923
rect 16715 13889 16724 13923
rect 16672 13880 16724 13889
rect 18604 13991 18656 14000
rect 18604 13957 18638 13991
rect 18638 13957 18656 13991
rect 18604 13948 18656 13957
rect 20168 14016 20220 14068
rect 20260 14016 20312 14068
rect 19984 13991 20036 14000
rect 19984 13957 19993 13991
rect 19993 13957 20027 13991
rect 20027 13957 20036 13991
rect 19984 13948 20036 13957
rect 20076 13991 20128 14000
rect 20076 13957 20085 13991
rect 20085 13957 20119 13991
rect 20119 13957 20128 13991
rect 20076 13948 20128 13957
rect 21640 14016 21692 14068
rect 22100 14016 22152 14068
rect 14556 13744 14608 13796
rect 14924 13744 14976 13796
rect 16580 13812 16632 13864
rect 21088 13880 21140 13932
rect 20812 13855 20864 13864
rect 20812 13821 20821 13855
rect 20821 13821 20855 13855
rect 20855 13821 20864 13855
rect 20812 13812 20864 13821
rect 21272 13812 21324 13864
rect 21732 13880 21784 13932
rect 23296 13880 23348 13932
rect 26424 14016 26476 14068
rect 27252 13948 27304 14000
rect 25780 13880 25832 13932
rect 26332 13923 26384 13932
rect 26332 13889 26341 13923
rect 26341 13889 26375 13923
rect 26375 13889 26384 13923
rect 26332 13880 26384 13889
rect 26700 13880 26752 13932
rect 31208 13923 31260 13932
rect 31208 13889 31217 13923
rect 31217 13889 31251 13923
rect 31251 13889 31260 13923
rect 31208 13880 31260 13889
rect 15384 13676 15436 13728
rect 15844 13676 15896 13728
rect 16028 13676 16080 13728
rect 22652 13744 22704 13796
rect 21732 13676 21784 13728
rect 29644 13812 29696 13864
rect 30104 13855 30156 13864
rect 30104 13821 30113 13855
rect 30113 13821 30147 13855
rect 30147 13821 30156 13855
rect 30104 13812 30156 13821
rect 31484 13855 31536 13864
rect 31484 13821 31493 13855
rect 31493 13821 31527 13855
rect 31527 13821 31536 13855
rect 31484 13812 31536 13821
rect 30012 13744 30064 13796
rect 25412 13719 25464 13728
rect 25412 13685 25421 13719
rect 25421 13685 25455 13719
rect 25455 13685 25464 13719
rect 25412 13676 25464 13685
rect 26148 13719 26200 13728
rect 26148 13685 26157 13719
rect 26157 13685 26191 13719
rect 26191 13685 26200 13719
rect 26148 13676 26200 13685
rect 27344 13719 27396 13728
rect 27344 13685 27353 13719
rect 27353 13685 27387 13719
rect 27387 13685 27396 13719
rect 27344 13676 27396 13685
rect 27436 13676 27488 13728
rect 27896 13676 27948 13728
rect 29368 13676 29420 13728
rect 4182 13574 4234 13626
rect 4246 13574 4298 13626
rect 4310 13574 4362 13626
rect 4374 13574 4426 13626
rect 4438 13574 4490 13626
rect 4502 13574 4554 13626
rect 10182 13574 10234 13626
rect 10246 13574 10298 13626
rect 10310 13574 10362 13626
rect 10374 13574 10426 13626
rect 10438 13574 10490 13626
rect 10502 13574 10554 13626
rect 16182 13574 16234 13626
rect 16246 13574 16298 13626
rect 16310 13574 16362 13626
rect 16374 13574 16426 13626
rect 16438 13574 16490 13626
rect 16502 13574 16554 13626
rect 22182 13574 22234 13626
rect 22246 13574 22298 13626
rect 22310 13574 22362 13626
rect 22374 13574 22426 13626
rect 22438 13574 22490 13626
rect 22502 13574 22554 13626
rect 28182 13574 28234 13626
rect 28246 13574 28298 13626
rect 28310 13574 28362 13626
rect 28374 13574 28426 13626
rect 28438 13574 28490 13626
rect 28502 13574 28554 13626
rect 3240 13472 3292 13524
rect 3792 13268 3844 13320
rect 14832 13472 14884 13524
rect 16212 13472 16264 13524
rect 18144 13472 18196 13524
rect 23296 13472 23348 13524
rect 14004 13404 14056 13456
rect 12532 13311 12584 13320
rect 12532 13277 12541 13311
rect 12541 13277 12575 13311
rect 12575 13277 12584 13311
rect 14096 13336 14148 13388
rect 14556 13379 14608 13388
rect 14556 13345 14565 13379
rect 14565 13345 14599 13379
rect 14599 13345 14608 13379
rect 14556 13336 14608 13345
rect 14648 13379 14700 13388
rect 14648 13345 14657 13379
rect 14657 13345 14691 13379
rect 14691 13345 14700 13379
rect 14648 13336 14700 13345
rect 22100 13404 22152 13456
rect 25780 13515 25832 13524
rect 25780 13481 25789 13515
rect 25789 13481 25823 13515
rect 25823 13481 25832 13515
rect 25780 13472 25832 13481
rect 27252 13515 27304 13524
rect 27252 13481 27261 13515
rect 27261 13481 27295 13515
rect 27295 13481 27304 13515
rect 27252 13472 27304 13481
rect 19708 13336 19760 13388
rect 12532 13268 12584 13277
rect 16028 13311 16080 13320
rect 16028 13277 16037 13311
rect 16037 13277 16071 13311
rect 16071 13277 16080 13311
rect 16028 13268 16080 13277
rect 16120 13311 16172 13320
rect 16120 13277 16129 13311
rect 16129 13277 16163 13311
rect 16163 13277 16172 13311
rect 16120 13268 16172 13277
rect 16212 13268 16264 13320
rect 16580 13311 16632 13320
rect 16580 13277 16589 13311
rect 16589 13277 16623 13311
rect 16623 13277 16632 13311
rect 16580 13268 16632 13277
rect 24032 13311 24084 13320
rect 24032 13277 24041 13311
rect 24041 13277 24075 13311
rect 24075 13277 24084 13311
rect 24032 13268 24084 13277
rect 26700 13268 26752 13320
rect 27896 13268 27948 13320
rect 28632 13268 28684 13320
rect 15660 13175 15712 13184
rect 15660 13141 15669 13175
rect 15669 13141 15703 13175
rect 15703 13141 15712 13175
rect 15660 13132 15712 13141
rect 16028 13132 16080 13184
rect 26148 13243 26200 13252
rect 26148 13209 26182 13243
rect 26182 13209 26200 13243
rect 26148 13200 26200 13209
rect 29368 13515 29420 13524
rect 29368 13481 29377 13515
rect 29377 13481 29411 13515
rect 29411 13481 29420 13515
rect 29368 13472 29420 13481
rect 29552 13472 29604 13524
rect 29920 13404 29972 13456
rect 30104 13311 30156 13320
rect 30104 13277 30112 13311
rect 30112 13277 30146 13311
rect 30146 13277 30156 13311
rect 30104 13268 30156 13277
rect 29828 13243 29880 13252
rect 29828 13209 29837 13243
rect 29837 13209 29871 13243
rect 29871 13209 29880 13243
rect 29828 13200 29880 13209
rect 30656 13200 30708 13252
rect 29736 13132 29788 13184
rect 30196 13132 30248 13184
rect 4922 13030 4974 13082
rect 4986 13030 5038 13082
rect 5050 13030 5102 13082
rect 5114 13030 5166 13082
rect 5178 13030 5230 13082
rect 5242 13030 5294 13082
rect 10922 13030 10974 13082
rect 10986 13030 11038 13082
rect 11050 13030 11102 13082
rect 11114 13030 11166 13082
rect 11178 13030 11230 13082
rect 11242 13030 11294 13082
rect 16922 13030 16974 13082
rect 16986 13030 17038 13082
rect 17050 13030 17102 13082
rect 17114 13030 17166 13082
rect 17178 13030 17230 13082
rect 17242 13030 17294 13082
rect 22922 13030 22974 13082
rect 22986 13030 23038 13082
rect 23050 13030 23102 13082
rect 23114 13030 23166 13082
rect 23178 13030 23230 13082
rect 23242 13030 23294 13082
rect 28922 13030 28974 13082
rect 28986 13030 29038 13082
rect 29050 13030 29102 13082
rect 29114 13030 29166 13082
rect 29178 13030 29230 13082
rect 29242 13030 29294 13082
rect 9772 12928 9824 12980
rect 14004 12928 14056 12980
rect 15936 12928 15988 12980
rect 22652 12928 22704 12980
rect 24032 12928 24084 12980
rect 25412 12928 25464 12980
rect 26332 12928 26384 12980
rect 27344 12971 27396 12980
rect 27344 12937 27353 12971
rect 27353 12937 27387 12971
rect 27387 12937 27396 12971
rect 27344 12928 27396 12937
rect 8300 12792 8352 12844
rect 9036 12860 9088 12912
rect 12900 12860 12952 12912
rect 13268 12860 13320 12912
rect 13452 12860 13504 12912
rect 8944 12767 8996 12776
rect 8944 12733 8953 12767
rect 8953 12733 8987 12767
rect 8987 12733 8996 12767
rect 8944 12724 8996 12733
rect 9680 12724 9732 12776
rect 12624 12792 12676 12844
rect 12808 12835 12860 12844
rect 12808 12801 12817 12835
rect 12817 12801 12851 12835
rect 12851 12801 12860 12835
rect 12808 12792 12860 12801
rect 13084 12835 13136 12844
rect 13084 12801 13093 12835
rect 13093 12801 13127 12835
rect 13127 12801 13136 12835
rect 13084 12792 13136 12801
rect 13820 12860 13872 12912
rect 10048 12656 10100 12708
rect 1492 12631 1544 12640
rect 1492 12597 1501 12631
rect 1501 12597 1535 12631
rect 1535 12597 1544 12631
rect 1492 12588 1544 12597
rect 14188 12792 14240 12844
rect 14372 12792 14424 12844
rect 20536 12835 20588 12844
rect 20536 12801 20545 12835
rect 20545 12801 20579 12835
rect 20579 12801 20588 12835
rect 20536 12792 20588 12801
rect 22928 12792 22980 12844
rect 25412 12792 25464 12844
rect 26700 12903 26752 12912
rect 26700 12869 26709 12903
rect 26709 12869 26743 12903
rect 26743 12869 26752 12903
rect 29368 12928 29420 12980
rect 29552 12928 29604 12980
rect 29828 12928 29880 12980
rect 26700 12860 26752 12869
rect 27436 12835 27488 12844
rect 27436 12801 27445 12835
rect 27445 12801 27479 12835
rect 27479 12801 27488 12835
rect 27436 12792 27488 12801
rect 21456 12724 21508 12776
rect 23848 12767 23900 12776
rect 23848 12733 23857 12767
rect 23857 12733 23891 12767
rect 23891 12733 23900 12767
rect 23848 12724 23900 12733
rect 25228 12724 25280 12776
rect 27068 12724 27120 12776
rect 27528 12767 27580 12776
rect 27528 12733 27537 12767
rect 27537 12733 27571 12767
rect 27571 12733 27580 12767
rect 27528 12724 27580 12733
rect 13544 12588 13596 12640
rect 22100 12588 22152 12640
rect 23296 12631 23348 12640
rect 23296 12597 23305 12631
rect 23305 12597 23339 12631
rect 23339 12597 23348 12631
rect 23296 12588 23348 12597
rect 28632 12835 28684 12844
rect 28632 12801 28641 12835
rect 28641 12801 28675 12835
rect 28675 12801 28684 12835
rect 28632 12792 28684 12801
rect 29552 12588 29604 12640
rect 30104 12631 30156 12640
rect 30104 12597 30113 12631
rect 30113 12597 30147 12631
rect 30147 12597 30156 12631
rect 30104 12588 30156 12597
rect 4182 12486 4234 12538
rect 4246 12486 4298 12538
rect 4310 12486 4362 12538
rect 4374 12486 4426 12538
rect 4438 12486 4490 12538
rect 4502 12486 4554 12538
rect 10182 12486 10234 12538
rect 10246 12486 10298 12538
rect 10310 12486 10362 12538
rect 10374 12486 10426 12538
rect 10438 12486 10490 12538
rect 10502 12486 10554 12538
rect 16182 12486 16234 12538
rect 16246 12486 16298 12538
rect 16310 12486 16362 12538
rect 16374 12486 16426 12538
rect 16438 12486 16490 12538
rect 16502 12486 16554 12538
rect 22182 12486 22234 12538
rect 22246 12486 22298 12538
rect 22310 12486 22362 12538
rect 22374 12486 22426 12538
rect 22438 12486 22490 12538
rect 22502 12486 22554 12538
rect 28182 12486 28234 12538
rect 28246 12486 28298 12538
rect 28310 12486 28362 12538
rect 28374 12486 28426 12538
rect 28438 12486 28490 12538
rect 28502 12486 28554 12538
rect 8944 12384 8996 12436
rect 22928 12427 22980 12436
rect 22928 12393 22937 12427
rect 22937 12393 22971 12427
rect 22971 12393 22980 12427
rect 22928 12384 22980 12393
rect 29552 12427 29604 12436
rect 29552 12393 29561 12427
rect 29561 12393 29595 12427
rect 29595 12393 29604 12427
rect 29552 12384 29604 12393
rect 5448 12316 5500 12368
rect 4160 12248 4212 12300
rect 4712 12248 4764 12300
rect 7196 12248 7248 12300
rect 4804 12180 4856 12232
rect 4712 12112 4764 12164
rect 7012 12223 7064 12232
rect 7012 12189 7021 12223
rect 7021 12189 7055 12223
rect 7055 12189 7064 12223
rect 7012 12180 7064 12189
rect 3976 12044 4028 12096
rect 4252 12087 4304 12096
rect 4252 12053 4261 12087
rect 4261 12053 4295 12087
rect 4295 12053 4304 12087
rect 4252 12044 4304 12053
rect 4436 12044 4488 12096
rect 6368 12087 6420 12096
rect 6368 12053 6377 12087
rect 6377 12053 6411 12087
rect 6411 12053 6420 12087
rect 6368 12044 6420 12053
rect 7104 12112 7156 12164
rect 9680 12316 9732 12368
rect 10048 12316 10100 12368
rect 9956 12291 10008 12300
rect 9956 12257 9965 12291
rect 9965 12257 9999 12291
rect 9999 12257 10008 12291
rect 9956 12248 10008 12257
rect 15292 12248 15344 12300
rect 15568 12248 15620 12300
rect 15844 12291 15896 12300
rect 15844 12257 15853 12291
rect 15853 12257 15887 12291
rect 15887 12257 15896 12291
rect 15844 12248 15896 12257
rect 8024 12223 8076 12232
rect 8024 12189 8033 12223
rect 8033 12189 8067 12223
rect 8067 12189 8076 12223
rect 8024 12180 8076 12189
rect 8668 12223 8720 12232
rect 8668 12189 8677 12223
rect 8677 12189 8711 12223
rect 8711 12189 8720 12223
rect 8668 12180 8720 12189
rect 6828 12087 6880 12096
rect 6828 12053 6837 12087
rect 6837 12053 6871 12087
rect 6871 12053 6880 12087
rect 6828 12044 6880 12053
rect 6920 12044 6972 12096
rect 7932 12044 7984 12096
rect 8484 12087 8536 12096
rect 8484 12053 8493 12087
rect 8493 12053 8527 12087
rect 8527 12053 8536 12087
rect 8484 12044 8536 12053
rect 9772 12223 9824 12232
rect 9772 12189 9781 12223
rect 9781 12189 9815 12223
rect 9815 12189 9824 12223
rect 9772 12180 9824 12189
rect 16120 12180 16172 12232
rect 21456 12291 21508 12300
rect 21456 12257 21465 12291
rect 21465 12257 21499 12291
rect 21499 12257 21508 12291
rect 21456 12248 21508 12257
rect 27528 12248 27580 12300
rect 30012 12291 30064 12300
rect 30012 12257 30021 12291
rect 30021 12257 30055 12291
rect 30055 12257 30064 12291
rect 30012 12248 30064 12257
rect 30196 12291 30248 12300
rect 30196 12257 30205 12291
rect 30205 12257 30239 12291
rect 30239 12257 30248 12291
rect 30196 12248 30248 12257
rect 23296 12223 23348 12232
rect 23296 12189 23305 12223
rect 23305 12189 23339 12223
rect 23339 12189 23348 12223
rect 23296 12180 23348 12189
rect 21272 12112 21324 12164
rect 10048 12044 10100 12096
rect 16028 12044 16080 12096
rect 19248 12087 19300 12096
rect 19248 12053 19257 12087
rect 19257 12053 19291 12087
rect 19291 12053 19300 12087
rect 19248 12044 19300 12053
rect 19708 12087 19760 12096
rect 19708 12053 19717 12087
rect 19717 12053 19751 12087
rect 19751 12053 19760 12087
rect 19708 12044 19760 12053
rect 21088 12044 21140 12096
rect 25412 12155 25464 12164
rect 25412 12121 25421 12155
rect 25421 12121 25455 12155
rect 25455 12121 25464 12155
rect 25412 12112 25464 12121
rect 26056 12112 26108 12164
rect 30104 12112 30156 12164
rect 22836 12087 22888 12096
rect 22836 12053 22845 12087
rect 22845 12053 22879 12087
rect 22879 12053 22888 12087
rect 22836 12044 22888 12053
rect 24676 12044 24728 12096
rect 4922 11942 4974 11994
rect 4986 11942 5038 11994
rect 5050 11942 5102 11994
rect 5114 11942 5166 11994
rect 5178 11942 5230 11994
rect 5242 11942 5294 11994
rect 10922 11942 10974 11994
rect 10986 11942 11038 11994
rect 11050 11942 11102 11994
rect 11114 11942 11166 11994
rect 11178 11942 11230 11994
rect 11242 11942 11294 11994
rect 16922 11942 16974 11994
rect 16986 11942 17038 11994
rect 17050 11942 17102 11994
rect 17114 11942 17166 11994
rect 17178 11942 17230 11994
rect 17242 11942 17294 11994
rect 22922 11942 22974 11994
rect 22986 11942 23038 11994
rect 23050 11942 23102 11994
rect 23114 11942 23166 11994
rect 23178 11942 23230 11994
rect 23242 11942 23294 11994
rect 28922 11942 28974 11994
rect 28986 11942 29038 11994
rect 29050 11942 29102 11994
rect 29114 11942 29166 11994
rect 29178 11942 29230 11994
rect 29242 11942 29294 11994
rect 3976 11883 4028 11892
rect 3976 11849 3985 11883
rect 3985 11849 4019 11883
rect 4019 11849 4028 11883
rect 3976 11840 4028 11849
rect 4252 11840 4304 11892
rect 4712 11840 4764 11892
rect 5080 11840 5132 11892
rect 5448 11840 5500 11892
rect 6368 11840 6420 11892
rect 6828 11840 6880 11892
rect 8024 11840 8076 11892
rect 16120 11840 16172 11892
rect 23848 11840 23900 11892
rect 2596 11747 2648 11756
rect 2596 11713 2605 11747
rect 2605 11713 2639 11747
rect 2639 11713 2648 11747
rect 2596 11704 2648 11713
rect 4436 11704 4488 11756
rect 4804 11704 4856 11756
rect 5080 11747 5132 11756
rect 5080 11713 5089 11747
rect 5089 11713 5123 11747
rect 5123 11713 5132 11747
rect 5080 11704 5132 11713
rect 5172 11747 5224 11756
rect 5172 11713 5181 11747
rect 5181 11713 5215 11747
rect 5215 11713 5224 11747
rect 5172 11704 5224 11713
rect 5356 11704 5408 11756
rect 6184 11704 6236 11756
rect 6368 11747 6420 11756
rect 6368 11713 6377 11747
rect 6377 11713 6411 11747
rect 6411 11713 6420 11747
rect 6368 11704 6420 11713
rect 3700 11636 3752 11688
rect 4160 11679 4212 11688
rect 4160 11645 4169 11679
rect 4169 11645 4203 11679
rect 4203 11645 4212 11679
rect 4160 11636 4212 11645
rect 5632 11679 5684 11688
rect 5632 11645 5641 11679
rect 5641 11645 5675 11679
rect 5675 11645 5684 11679
rect 7932 11704 7984 11756
rect 5632 11636 5684 11645
rect 7380 11636 7432 11688
rect 9864 11704 9916 11756
rect 14188 11704 14240 11756
rect 15936 11704 15988 11756
rect 17960 11747 18012 11756
rect 17960 11713 17994 11747
rect 17994 11713 18012 11747
rect 17960 11704 18012 11713
rect 8944 11636 8996 11688
rect 14004 11636 14056 11688
rect 19432 11747 19484 11756
rect 19432 11713 19466 11747
rect 19466 11713 19484 11747
rect 19432 11704 19484 11713
rect 20720 11772 20772 11824
rect 21640 11772 21692 11824
rect 22100 11815 22152 11824
rect 22100 11781 22134 11815
rect 22134 11781 22152 11815
rect 22100 11772 22152 11781
rect 22284 11772 22336 11824
rect 26516 11815 26568 11824
rect 26516 11781 26525 11815
rect 26525 11781 26559 11815
rect 26559 11781 26568 11815
rect 26516 11772 26568 11781
rect 22836 11704 22888 11756
rect 23480 11704 23532 11756
rect 25780 11747 25832 11756
rect 25780 11713 25789 11747
rect 25789 11713 25823 11747
rect 25823 11713 25832 11747
rect 25780 11704 25832 11713
rect 26332 11747 26384 11756
rect 26332 11713 26341 11747
rect 26341 11713 26375 11747
rect 26375 11713 26384 11747
rect 26332 11704 26384 11713
rect 6736 11500 6788 11552
rect 13084 11500 13136 11552
rect 14096 11500 14148 11552
rect 26700 11747 26752 11756
rect 26700 11713 26709 11747
rect 26709 11713 26743 11747
rect 26743 11713 26752 11747
rect 26700 11704 26752 11713
rect 28080 11636 28132 11688
rect 18972 11500 19024 11552
rect 20352 11500 20404 11552
rect 21088 11500 21140 11552
rect 21180 11500 21232 11552
rect 23388 11500 23440 11552
rect 25596 11543 25648 11552
rect 25596 11509 25605 11543
rect 25605 11509 25639 11543
rect 25639 11509 25648 11543
rect 25596 11500 25648 11509
rect 26424 11500 26476 11552
rect 26516 11500 26568 11552
rect 4182 11398 4234 11450
rect 4246 11398 4298 11450
rect 4310 11398 4362 11450
rect 4374 11398 4426 11450
rect 4438 11398 4490 11450
rect 4502 11398 4554 11450
rect 10182 11398 10234 11450
rect 10246 11398 10298 11450
rect 10310 11398 10362 11450
rect 10374 11398 10426 11450
rect 10438 11398 10490 11450
rect 10502 11398 10554 11450
rect 16182 11398 16234 11450
rect 16246 11398 16298 11450
rect 16310 11398 16362 11450
rect 16374 11398 16426 11450
rect 16438 11398 16490 11450
rect 16502 11398 16554 11450
rect 22182 11398 22234 11450
rect 22246 11398 22298 11450
rect 22310 11398 22362 11450
rect 22374 11398 22426 11450
rect 22438 11398 22490 11450
rect 22502 11398 22554 11450
rect 28182 11398 28234 11450
rect 28246 11398 28298 11450
rect 28310 11398 28362 11450
rect 28374 11398 28426 11450
rect 28438 11398 28490 11450
rect 28502 11398 28554 11450
rect 2596 11296 2648 11348
rect 3700 11296 3752 11348
rect 5632 11296 5684 11348
rect 6184 11296 6236 11348
rect 7380 11296 7432 11348
rect 14096 11296 14148 11348
rect 16028 11296 16080 11348
rect 17960 11296 18012 11348
rect 19432 11296 19484 11348
rect 21272 11296 21324 11348
rect 22836 11296 22888 11348
rect 25228 11296 25280 11348
rect 26700 11296 26752 11348
rect 28080 11339 28132 11348
rect 28080 11305 28089 11339
rect 28089 11305 28123 11339
rect 28123 11305 28132 11339
rect 28080 11296 28132 11305
rect 4068 11160 4120 11212
rect 8576 11228 8628 11280
rect 5908 11160 5960 11212
rect 5172 11135 5224 11144
rect 5172 11101 5181 11135
rect 5181 11101 5215 11135
rect 5215 11101 5224 11135
rect 5172 11092 5224 11101
rect 6368 11092 6420 11144
rect 7104 11092 7156 11144
rect 11336 11160 11388 11212
rect 13728 11160 13780 11212
rect 16120 11228 16172 11280
rect 9036 11135 9088 11144
rect 9036 11101 9045 11135
rect 9045 11101 9079 11135
rect 9079 11101 9088 11135
rect 9036 11092 9088 11101
rect 11520 11092 11572 11144
rect 12992 11135 13044 11144
rect 8484 11024 8536 11076
rect 9864 11067 9916 11076
rect 9864 11033 9873 11067
rect 9873 11033 9907 11067
rect 9907 11033 9916 11067
rect 12992 11101 13001 11135
rect 13001 11101 13035 11135
rect 13035 11101 13044 11135
rect 14096 11135 14148 11144
rect 12992 11092 13044 11101
rect 9864 11024 9916 11033
rect 13728 11067 13780 11076
rect 13728 11033 13737 11067
rect 13737 11033 13771 11067
rect 13771 11033 13780 11067
rect 13728 11024 13780 11033
rect 14096 11101 14105 11135
rect 14105 11101 14139 11135
rect 14139 11101 14148 11135
rect 14096 11092 14148 11101
rect 20352 11160 20404 11212
rect 19248 11092 19300 11144
rect 22100 11160 22152 11212
rect 21088 11067 21140 11076
rect 21088 11033 21097 11067
rect 21097 11033 21131 11067
rect 21131 11033 21140 11067
rect 21088 11024 21140 11033
rect 21180 11067 21232 11076
rect 21180 11033 21189 11067
rect 21189 11033 21223 11067
rect 21223 11033 21232 11067
rect 21180 11024 21232 11033
rect 22744 11092 22796 11144
rect 23112 11067 23164 11076
rect 23112 11033 23121 11067
rect 23121 11033 23155 11067
rect 23155 11033 23164 11067
rect 23112 11024 23164 11033
rect 23480 11092 23532 11144
rect 23848 11092 23900 11144
rect 25228 11135 25280 11144
rect 25228 11101 25237 11135
rect 25237 11101 25271 11135
rect 25271 11101 25280 11135
rect 25228 11092 25280 11101
rect 26056 11092 26108 11144
rect 25596 11024 25648 11076
rect 26792 11024 26844 11076
rect 9956 10999 10008 11008
rect 9956 10965 9965 10999
rect 9965 10965 9999 10999
rect 9999 10965 10008 10999
rect 9956 10956 10008 10965
rect 10692 10999 10744 11008
rect 10692 10965 10701 10999
rect 10701 10965 10735 10999
rect 10735 10965 10744 10999
rect 10692 10956 10744 10965
rect 12348 10999 12400 11008
rect 12348 10965 12357 10999
rect 12357 10965 12391 10999
rect 12391 10965 12400 10999
rect 12348 10956 12400 10965
rect 13820 10956 13872 11008
rect 15476 10999 15528 11008
rect 15476 10965 15485 10999
rect 15485 10965 15519 10999
rect 15519 10965 15528 10999
rect 15476 10956 15528 10965
rect 15568 10999 15620 11008
rect 15568 10965 15577 10999
rect 15577 10965 15611 10999
rect 15611 10965 15620 10999
rect 15568 10956 15620 10965
rect 19432 10956 19484 11008
rect 19708 10999 19760 11008
rect 19708 10965 19717 10999
rect 19717 10965 19751 10999
rect 19751 10965 19760 10999
rect 19708 10956 19760 10965
rect 20812 10999 20864 11008
rect 20812 10965 20821 10999
rect 20821 10965 20855 10999
rect 20855 10965 20864 10999
rect 20812 10956 20864 10965
rect 24676 10956 24728 11008
rect 28172 10999 28224 11008
rect 28172 10965 28181 10999
rect 28181 10965 28215 10999
rect 28215 10965 28224 10999
rect 28172 10956 28224 10965
rect 4922 10854 4974 10906
rect 4986 10854 5038 10906
rect 5050 10854 5102 10906
rect 5114 10854 5166 10906
rect 5178 10854 5230 10906
rect 5242 10854 5294 10906
rect 10922 10854 10974 10906
rect 10986 10854 11038 10906
rect 11050 10854 11102 10906
rect 11114 10854 11166 10906
rect 11178 10854 11230 10906
rect 11242 10854 11294 10906
rect 16922 10854 16974 10906
rect 16986 10854 17038 10906
rect 17050 10854 17102 10906
rect 17114 10854 17166 10906
rect 17178 10854 17230 10906
rect 17242 10854 17294 10906
rect 22922 10854 22974 10906
rect 22986 10854 23038 10906
rect 23050 10854 23102 10906
rect 23114 10854 23166 10906
rect 23178 10854 23230 10906
rect 23242 10854 23294 10906
rect 28922 10854 28974 10906
rect 28986 10854 29038 10906
rect 29050 10854 29102 10906
rect 29114 10854 29166 10906
rect 29178 10854 29230 10906
rect 29242 10854 29294 10906
rect 4712 10684 4764 10736
rect 2596 10616 2648 10668
rect 5172 10616 5224 10668
rect 2504 10591 2556 10600
rect 2504 10557 2513 10591
rect 2513 10557 2547 10591
rect 2547 10557 2556 10591
rect 2504 10548 2556 10557
rect 4620 10591 4672 10600
rect 4620 10557 4629 10591
rect 4629 10557 4663 10591
rect 4663 10557 4672 10591
rect 4620 10548 4672 10557
rect 5632 10616 5684 10668
rect 6920 10795 6972 10804
rect 6920 10761 6929 10795
rect 6929 10761 6963 10795
rect 6963 10761 6972 10795
rect 6920 10752 6972 10761
rect 7012 10752 7064 10804
rect 8392 10752 8444 10804
rect 8576 10752 8628 10804
rect 8668 10752 8720 10804
rect 9956 10752 10008 10804
rect 11336 10795 11388 10804
rect 11336 10761 11345 10795
rect 11345 10761 11379 10795
rect 11379 10761 11388 10795
rect 11336 10752 11388 10761
rect 11520 10795 11572 10804
rect 11520 10761 11529 10795
rect 11529 10761 11563 10795
rect 11563 10761 11572 10795
rect 11520 10752 11572 10761
rect 12348 10752 12400 10804
rect 14188 10795 14240 10804
rect 14188 10761 14197 10795
rect 14197 10761 14231 10795
rect 14231 10761 14240 10795
rect 14188 10752 14240 10761
rect 15568 10752 15620 10804
rect 25780 10752 25832 10804
rect 26516 10752 26568 10804
rect 26792 10752 26844 10804
rect 28172 10752 28224 10804
rect 7196 10684 7248 10736
rect 6184 10548 6236 10600
rect 3976 10455 4028 10464
rect 3976 10421 3985 10455
rect 3985 10421 4019 10455
rect 4019 10421 4028 10455
rect 3976 10412 4028 10421
rect 4068 10412 4120 10464
rect 6736 10548 6788 10600
rect 10692 10684 10744 10736
rect 10876 10684 10928 10736
rect 11612 10684 11664 10736
rect 13820 10727 13872 10736
rect 13820 10693 13829 10727
rect 13829 10693 13863 10727
rect 13863 10693 13872 10727
rect 13820 10684 13872 10693
rect 24400 10684 24452 10736
rect 29368 10752 29420 10804
rect 29736 10752 29788 10804
rect 15108 10616 15160 10668
rect 19524 10616 19576 10668
rect 20260 10616 20312 10668
rect 20352 10659 20404 10668
rect 20352 10625 20361 10659
rect 20361 10625 20395 10659
rect 20395 10625 20404 10659
rect 20352 10616 20404 10625
rect 8576 10548 8628 10600
rect 8760 10412 8812 10464
rect 8852 10455 8904 10464
rect 8852 10421 8861 10455
rect 8861 10421 8895 10455
rect 8895 10421 8904 10455
rect 8852 10412 8904 10421
rect 9036 10480 9088 10532
rect 12164 10591 12216 10600
rect 12164 10557 12173 10591
rect 12173 10557 12207 10591
rect 12207 10557 12216 10591
rect 12164 10548 12216 10557
rect 15292 10548 15344 10600
rect 19708 10591 19760 10600
rect 19708 10557 19717 10591
rect 19717 10557 19751 10591
rect 19751 10557 19760 10591
rect 19708 10548 19760 10557
rect 25320 10548 25372 10600
rect 14096 10412 14148 10464
rect 14832 10412 14884 10464
rect 20076 10455 20128 10464
rect 20076 10421 20085 10455
rect 20085 10421 20119 10455
rect 20119 10421 20128 10455
rect 20076 10412 20128 10421
rect 20168 10455 20220 10464
rect 20168 10421 20177 10455
rect 20177 10421 20211 10455
rect 20211 10421 20220 10455
rect 20168 10412 20220 10421
rect 20812 10412 20864 10464
rect 27436 10591 27488 10600
rect 27436 10557 27445 10591
rect 27445 10557 27479 10591
rect 27479 10557 27488 10591
rect 27436 10548 27488 10557
rect 27528 10591 27580 10600
rect 27528 10557 27537 10591
rect 27537 10557 27571 10591
rect 27571 10557 27580 10591
rect 27528 10548 27580 10557
rect 30196 10548 30248 10600
rect 29000 10412 29052 10464
rect 4182 10310 4234 10362
rect 4246 10310 4298 10362
rect 4310 10310 4362 10362
rect 4374 10310 4426 10362
rect 4438 10310 4490 10362
rect 4502 10310 4554 10362
rect 10182 10310 10234 10362
rect 10246 10310 10298 10362
rect 10310 10310 10362 10362
rect 10374 10310 10426 10362
rect 10438 10310 10490 10362
rect 10502 10310 10554 10362
rect 16182 10310 16234 10362
rect 16246 10310 16298 10362
rect 16310 10310 16362 10362
rect 16374 10310 16426 10362
rect 16438 10310 16490 10362
rect 16502 10310 16554 10362
rect 22182 10310 22234 10362
rect 22246 10310 22298 10362
rect 22310 10310 22362 10362
rect 22374 10310 22426 10362
rect 22438 10310 22490 10362
rect 22502 10310 22554 10362
rect 28182 10310 28234 10362
rect 28246 10310 28298 10362
rect 28310 10310 28362 10362
rect 28374 10310 28426 10362
rect 28438 10310 28490 10362
rect 28502 10310 28554 10362
rect 2596 10251 2648 10260
rect 2596 10217 2605 10251
rect 2605 10217 2639 10251
rect 2639 10217 2648 10251
rect 2596 10208 2648 10217
rect 3976 10208 4028 10260
rect 8484 10208 8536 10260
rect 8852 10208 8904 10260
rect 10048 10208 10100 10260
rect 4068 10072 4120 10124
rect 20076 10208 20128 10260
rect 20260 10208 20312 10260
rect 23756 10208 23808 10260
rect 29920 10208 29972 10260
rect 4712 10004 4764 10056
rect 5172 10047 5224 10056
rect 5172 10013 5181 10047
rect 5181 10013 5215 10047
rect 5215 10013 5224 10047
rect 5172 10004 5224 10013
rect 8392 10004 8444 10056
rect 9864 9936 9916 9988
rect 11336 10004 11388 10056
rect 12900 10004 12952 10056
rect 13084 10004 13136 10056
rect 14096 10047 14148 10056
rect 14096 10013 14105 10047
rect 14105 10013 14139 10047
rect 14139 10013 14148 10047
rect 14096 10004 14148 10013
rect 11796 9936 11848 9988
rect 15476 10072 15528 10124
rect 25044 10140 25096 10192
rect 14832 10047 14884 10056
rect 14832 10013 14841 10047
rect 14841 10013 14875 10047
rect 14875 10013 14884 10047
rect 14832 10004 14884 10013
rect 20260 10004 20312 10056
rect 24584 10072 24636 10124
rect 14924 9936 14976 9988
rect 3792 9911 3844 9920
rect 3792 9877 3801 9911
rect 3801 9877 3835 9911
rect 3835 9877 3844 9911
rect 3792 9868 3844 9877
rect 4528 9868 4580 9920
rect 7932 9911 7984 9920
rect 7932 9877 7941 9911
rect 7941 9877 7975 9911
rect 7975 9877 7984 9911
rect 7932 9868 7984 9877
rect 8576 9868 8628 9920
rect 11520 9911 11572 9920
rect 11520 9877 11529 9911
rect 11529 9877 11563 9911
rect 11563 9877 11572 9911
rect 11520 9868 11572 9877
rect 14648 9911 14700 9920
rect 14648 9877 14657 9911
rect 14657 9877 14691 9911
rect 14691 9877 14700 9911
rect 14648 9868 14700 9877
rect 19340 9911 19392 9920
rect 19340 9877 19349 9911
rect 19349 9877 19383 9911
rect 19383 9877 19392 9911
rect 19340 9868 19392 9877
rect 19432 9868 19484 9920
rect 21180 9979 21232 9988
rect 21180 9945 21189 9979
rect 21189 9945 21223 9979
rect 21223 9945 21232 9979
rect 21180 9936 21232 9945
rect 21272 9979 21324 9988
rect 21272 9945 21281 9979
rect 21281 9945 21315 9979
rect 21315 9945 21324 9979
rect 21272 9936 21324 9945
rect 24308 9936 24360 9988
rect 23756 9868 23808 9920
rect 24492 10004 24544 10056
rect 26056 10004 26108 10056
rect 30104 10115 30156 10124
rect 30104 10081 30113 10115
rect 30113 10081 30147 10115
rect 30147 10081 30156 10115
rect 30104 10072 30156 10081
rect 30196 10072 30248 10124
rect 29736 10004 29788 10056
rect 30656 9979 30708 9988
rect 30656 9945 30665 9979
rect 30665 9945 30699 9979
rect 30699 9945 30708 9979
rect 30656 9936 30708 9945
rect 30748 9979 30800 9988
rect 30748 9945 30757 9979
rect 30757 9945 30791 9979
rect 30791 9945 30800 9979
rect 30748 9936 30800 9945
rect 24676 9868 24728 9920
rect 29460 9868 29512 9920
rect 30012 9911 30064 9920
rect 30012 9877 30021 9911
rect 30021 9877 30055 9911
rect 30055 9877 30064 9911
rect 30012 9868 30064 9877
rect 30472 9868 30524 9920
rect 31024 9911 31076 9920
rect 31024 9877 31033 9911
rect 31033 9877 31067 9911
rect 31067 9877 31076 9911
rect 31024 9868 31076 9877
rect 4922 9766 4974 9818
rect 4986 9766 5038 9818
rect 5050 9766 5102 9818
rect 5114 9766 5166 9818
rect 5178 9766 5230 9818
rect 5242 9766 5294 9818
rect 10922 9766 10974 9818
rect 10986 9766 11038 9818
rect 11050 9766 11102 9818
rect 11114 9766 11166 9818
rect 11178 9766 11230 9818
rect 11242 9766 11294 9818
rect 16922 9766 16974 9818
rect 16986 9766 17038 9818
rect 17050 9766 17102 9818
rect 17114 9766 17166 9818
rect 17178 9766 17230 9818
rect 17242 9766 17294 9818
rect 22922 9766 22974 9818
rect 22986 9766 23038 9818
rect 23050 9766 23102 9818
rect 23114 9766 23166 9818
rect 23178 9766 23230 9818
rect 23242 9766 23294 9818
rect 28922 9766 28974 9818
rect 28986 9766 29038 9818
rect 29050 9766 29102 9818
rect 29114 9766 29166 9818
rect 29178 9766 29230 9818
rect 29242 9766 29294 9818
rect 7196 9664 7248 9716
rect 8392 9707 8444 9716
rect 8392 9673 8401 9707
rect 8401 9673 8435 9707
rect 8435 9673 8444 9707
rect 8392 9664 8444 9673
rect 11244 9664 11296 9716
rect 12900 9707 12952 9716
rect 12900 9673 12909 9707
rect 12909 9673 12943 9707
rect 12943 9673 12952 9707
rect 12900 9664 12952 9673
rect 2504 9571 2556 9580
rect 2504 9537 2513 9571
rect 2513 9537 2547 9571
rect 2547 9537 2556 9571
rect 2504 9528 2556 9537
rect 2780 9571 2832 9580
rect 2780 9537 2814 9571
rect 2814 9537 2832 9571
rect 2780 9528 2832 9537
rect 7288 9571 7340 9580
rect 7288 9537 7322 9571
rect 7322 9537 7340 9571
rect 7288 9528 7340 9537
rect 11152 9571 11204 9580
rect 11152 9537 11161 9571
rect 11161 9537 11195 9571
rect 11195 9537 11204 9571
rect 11152 9528 11204 9537
rect 11612 9528 11664 9580
rect 14648 9596 14700 9648
rect 15752 9596 15804 9648
rect 20260 9707 20312 9716
rect 20260 9673 20269 9707
rect 20269 9673 20303 9707
rect 20303 9673 20312 9707
rect 20260 9664 20312 9673
rect 20352 9707 20404 9716
rect 20352 9673 20361 9707
rect 20361 9673 20395 9707
rect 20395 9673 20404 9707
rect 20352 9664 20404 9673
rect 21272 9664 21324 9716
rect 23664 9664 23716 9716
rect 25136 9639 25188 9648
rect 13820 9528 13872 9580
rect 6920 9460 6972 9512
rect 4712 9392 4764 9444
rect 12992 9367 13044 9376
rect 12992 9333 13001 9367
rect 13001 9333 13035 9367
rect 13035 9333 13044 9367
rect 12992 9324 13044 9333
rect 15384 9367 15436 9376
rect 15384 9333 15393 9367
rect 15393 9333 15427 9367
rect 15427 9333 15436 9367
rect 15384 9324 15436 9333
rect 15752 9324 15804 9376
rect 18972 9528 19024 9580
rect 19432 9528 19484 9580
rect 20720 9571 20772 9580
rect 20720 9537 20729 9571
rect 20729 9537 20763 9571
rect 20763 9537 20772 9571
rect 20720 9528 20772 9537
rect 23112 9571 23164 9580
rect 23112 9537 23121 9571
rect 23121 9537 23155 9571
rect 23155 9537 23164 9571
rect 23112 9528 23164 9537
rect 25136 9605 25148 9639
rect 25148 9605 25188 9639
rect 25136 9596 25188 9605
rect 28080 9596 28132 9648
rect 30012 9664 30064 9716
rect 30196 9707 30248 9716
rect 30196 9673 30205 9707
rect 30205 9673 30239 9707
rect 30239 9673 30248 9707
rect 30196 9664 30248 9673
rect 30472 9707 30524 9716
rect 30472 9673 30481 9707
rect 30481 9673 30515 9707
rect 30515 9673 30524 9707
rect 30472 9664 30524 9673
rect 28816 9596 28868 9648
rect 29092 9639 29144 9648
rect 29092 9605 29126 9639
rect 29126 9605 29144 9639
rect 29092 9596 29144 9605
rect 29644 9596 29696 9648
rect 24952 9528 25004 9580
rect 25688 9528 25740 9580
rect 30748 9528 30800 9580
rect 19248 9324 19300 9376
rect 28816 9503 28868 9512
rect 28816 9469 28832 9503
rect 28832 9469 28866 9503
rect 28866 9469 28868 9503
rect 28816 9460 28868 9469
rect 24492 9324 24544 9376
rect 24768 9367 24820 9376
rect 24768 9333 24777 9367
rect 24777 9333 24811 9367
rect 24811 9333 24820 9367
rect 24768 9324 24820 9333
rect 26056 9324 26108 9376
rect 28724 9367 28776 9376
rect 28724 9333 28733 9367
rect 28733 9333 28767 9367
rect 28767 9333 28776 9367
rect 28724 9324 28776 9333
rect 4182 9222 4234 9274
rect 4246 9222 4298 9274
rect 4310 9222 4362 9274
rect 4374 9222 4426 9274
rect 4438 9222 4490 9274
rect 4502 9222 4554 9274
rect 10182 9222 10234 9274
rect 10246 9222 10298 9274
rect 10310 9222 10362 9274
rect 10374 9222 10426 9274
rect 10438 9222 10490 9274
rect 10502 9222 10554 9274
rect 16182 9222 16234 9274
rect 16246 9222 16298 9274
rect 16310 9222 16362 9274
rect 16374 9222 16426 9274
rect 16438 9222 16490 9274
rect 16502 9222 16554 9274
rect 22182 9222 22234 9274
rect 22246 9222 22298 9274
rect 22310 9222 22362 9274
rect 22374 9222 22426 9274
rect 22438 9222 22490 9274
rect 22502 9222 22554 9274
rect 28182 9222 28234 9274
rect 28246 9222 28298 9274
rect 28310 9222 28362 9274
rect 28374 9222 28426 9274
rect 28438 9222 28490 9274
rect 28502 9222 28554 9274
rect 2780 9120 2832 9172
rect 7288 9120 7340 9172
rect 11152 9120 11204 9172
rect 14832 9120 14884 9172
rect 15384 9120 15436 9172
rect 18512 9120 18564 9172
rect 19708 9120 19760 9172
rect 20720 9120 20772 9172
rect 22836 9163 22888 9172
rect 22836 9129 22845 9163
rect 22845 9129 22879 9163
rect 22879 9129 22888 9163
rect 22836 9120 22888 9129
rect 23112 9120 23164 9172
rect 8760 9052 8812 9104
rect 11336 9052 11388 9104
rect 12164 8984 12216 9036
rect 15016 8984 15068 9036
rect 3792 8916 3844 8968
rect 7932 8916 7984 8968
rect 9772 8916 9824 8968
rect 10692 8848 10744 8900
rect 11520 8916 11572 8968
rect 12992 8916 13044 8968
rect 19340 9052 19392 9104
rect 8576 8780 8628 8832
rect 10324 8780 10376 8832
rect 10784 8823 10836 8832
rect 10784 8789 10793 8823
rect 10793 8789 10827 8823
rect 10827 8789 10836 8823
rect 10784 8780 10836 8789
rect 12440 8780 12492 8832
rect 13820 8780 13872 8832
rect 14372 8780 14424 8832
rect 15108 8780 15160 8832
rect 16488 8780 16540 8832
rect 17684 8780 17736 8832
rect 18052 8848 18104 8900
rect 18512 8959 18564 8968
rect 18512 8925 18521 8959
rect 18521 8925 18555 8959
rect 18555 8925 18564 8959
rect 18512 8916 18564 8925
rect 18696 8891 18748 8900
rect 18696 8857 18705 8891
rect 18705 8857 18739 8891
rect 18739 8857 18748 8891
rect 18696 8848 18748 8857
rect 18972 8916 19024 8968
rect 19892 8916 19944 8968
rect 20168 8916 20220 8968
rect 19432 8848 19484 8900
rect 26056 9120 26108 9172
rect 26424 9163 26476 9172
rect 26424 9129 26433 9163
rect 26433 9129 26467 9163
rect 26467 9129 26476 9163
rect 26424 9120 26476 9129
rect 28724 9120 28776 9172
rect 29092 9120 29144 9172
rect 30748 9120 30800 9172
rect 21180 8984 21232 9036
rect 21824 8984 21876 9036
rect 22652 8984 22704 9036
rect 22744 8959 22796 8968
rect 22744 8925 22753 8959
rect 22753 8925 22787 8959
rect 22787 8925 22796 8959
rect 22744 8916 22796 8925
rect 23756 8959 23808 8968
rect 22652 8848 22704 8900
rect 22100 8780 22152 8832
rect 22836 8780 22888 8832
rect 23756 8925 23760 8959
rect 23760 8925 23794 8959
rect 23794 8925 23808 8959
rect 23756 8916 23808 8925
rect 24768 9052 24820 9104
rect 24400 8916 24452 8968
rect 24584 8916 24636 8968
rect 25688 8984 25740 9036
rect 26608 8959 26660 8968
rect 26608 8925 26617 8959
rect 26617 8925 26651 8959
rect 26651 8925 26660 8959
rect 26608 8916 26660 8925
rect 28816 8984 28868 9036
rect 23664 8780 23716 8832
rect 26424 8891 26476 8900
rect 26424 8857 26433 8891
rect 26433 8857 26467 8891
rect 26467 8857 26476 8891
rect 26424 8848 26476 8857
rect 29460 8916 29512 8968
rect 31024 8916 31076 8968
rect 24860 8823 24912 8832
rect 24860 8789 24869 8823
rect 24869 8789 24903 8823
rect 24903 8789 24912 8823
rect 24860 8780 24912 8789
rect 26884 8823 26936 8832
rect 26884 8789 26893 8823
rect 26893 8789 26927 8823
rect 26927 8789 26936 8823
rect 26884 8780 26936 8789
rect 4922 8678 4974 8730
rect 4986 8678 5038 8730
rect 5050 8678 5102 8730
rect 5114 8678 5166 8730
rect 5178 8678 5230 8730
rect 5242 8678 5294 8730
rect 10922 8678 10974 8730
rect 10986 8678 11038 8730
rect 11050 8678 11102 8730
rect 11114 8678 11166 8730
rect 11178 8678 11230 8730
rect 11242 8678 11294 8730
rect 16922 8678 16974 8730
rect 16986 8678 17038 8730
rect 17050 8678 17102 8730
rect 17114 8678 17166 8730
rect 17178 8678 17230 8730
rect 17242 8678 17294 8730
rect 22922 8678 22974 8730
rect 22986 8678 23038 8730
rect 23050 8678 23102 8730
rect 23114 8678 23166 8730
rect 23178 8678 23230 8730
rect 23242 8678 23294 8730
rect 28922 8678 28974 8730
rect 28986 8678 29038 8730
rect 29050 8678 29102 8730
rect 29114 8678 29166 8730
rect 29178 8678 29230 8730
rect 29242 8678 29294 8730
rect 9864 8619 9916 8628
rect 9864 8585 9873 8619
rect 9873 8585 9907 8619
rect 9907 8585 9916 8619
rect 9864 8576 9916 8585
rect 10784 8576 10836 8628
rect 6000 8483 6052 8492
rect 6000 8449 6009 8483
rect 6009 8449 6043 8483
rect 6043 8449 6052 8483
rect 6000 8440 6052 8449
rect 6644 8372 6696 8424
rect 5816 8347 5868 8356
rect 5816 8313 5825 8347
rect 5825 8313 5859 8347
rect 5859 8313 5868 8347
rect 5816 8304 5868 8313
rect 8392 8483 8444 8492
rect 8392 8449 8401 8483
rect 8401 8449 8435 8483
rect 8435 8449 8444 8483
rect 8392 8440 8444 8449
rect 8944 8440 8996 8492
rect 9220 8483 9272 8492
rect 9220 8449 9229 8483
rect 9229 8449 9263 8483
rect 9263 8449 9272 8483
rect 9220 8440 9272 8449
rect 9956 8508 10008 8560
rect 13820 8576 13872 8628
rect 14004 8576 14056 8628
rect 15752 8576 15804 8628
rect 16488 8576 16540 8628
rect 18052 8619 18104 8628
rect 18052 8585 18061 8619
rect 18061 8585 18095 8619
rect 18095 8585 18104 8619
rect 18052 8576 18104 8585
rect 9680 8440 9732 8492
rect 8300 8304 8352 8356
rect 8484 8304 8536 8356
rect 9312 8304 9364 8356
rect 10048 8304 10100 8356
rect 10324 8372 10376 8424
rect 12440 8440 12492 8492
rect 13728 8440 13780 8492
rect 14096 8483 14148 8492
rect 14096 8449 14103 8483
rect 14103 8449 14148 8483
rect 14096 8440 14148 8449
rect 10784 8415 10836 8424
rect 10784 8381 10793 8415
rect 10793 8381 10827 8415
rect 10827 8381 10836 8415
rect 10784 8372 10836 8381
rect 15476 8508 15528 8560
rect 14372 8483 14424 8492
rect 14372 8449 14386 8483
rect 14386 8449 14420 8483
rect 14420 8449 14424 8483
rect 14372 8440 14424 8449
rect 14556 8440 14608 8492
rect 14832 8483 14884 8492
rect 14832 8449 14841 8483
rect 14841 8449 14875 8483
rect 14875 8449 14884 8483
rect 14832 8440 14884 8449
rect 14924 8483 14976 8492
rect 14924 8449 14933 8483
rect 14933 8449 14967 8483
rect 14967 8449 14976 8483
rect 14924 8440 14976 8449
rect 16672 8483 16724 8492
rect 16672 8449 16681 8483
rect 16681 8449 16715 8483
rect 16715 8449 16724 8483
rect 16672 8440 16724 8449
rect 19156 8576 19208 8628
rect 19432 8576 19484 8628
rect 20444 8576 20496 8628
rect 18696 8508 18748 8560
rect 19984 8508 20036 8560
rect 22100 8551 22152 8560
rect 22100 8517 22109 8551
rect 22109 8517 22143 8551
rect 22143 8517 22152 8551
rect 22100 8508 22152 8517
rect 6552 8236 6604 8288
rect 8668 8279 8720 8288
rect 8668 8245 8677 8279
rect 8677 8245 8711 8279
rect 8711 8245 8720 8279
rect 8668 8236 8720 8245
rect 9864 8236 9916 8288
rect 10784 8236 10836 8288
rect 16856 8236 16908 8288
rect 17316 8236 17368 8288
rect 19432 8372 19484 8424
rect 22192 8483 22244 8492
rect 22192 8449 22201 8483
rect 22201 8449 22235 8483
rect 22235 8449 22244 8483
rect 22192 8440 22244 8449
rect 22744 8576 22796 8628
rect 26608 8576 26660 8628
rect 22836 8508 22888 8560
rect 27344 8576 27396 8628
rect 18512 8304 18564 8356
rect 23388 8372 23440 8424
rect 27068 8372 27120 8424
rect 29368 8440 29420 8492
rect 22744 8304 22796 8356
rect 24676 8236 24728 8288
rect 28080 8304 28132 8356
rect 27436 8236 27488 8288
rect 27804 8279 27856 8288
rect 27804 8245 27813 8279
rect 27813 8245 27847 8279
rect 27847 8245 27856 8279
rect 27804 8236 27856 8245
rect 4182 8134 4234 8186
rect 4246 8134 4298 8186
rect 4310 8134 4362 8186
rect 4374 8134 4426 8186
rect 4438 8134 4490 8186
rect 4502 8134 4554 8186
rect 10182 8134 10234 8186
rect 10246 8134 10298 8186
rect 10310 8134 10362 8186
rect 10374 8134 10426 8186
rect 10438 8134 10490 8186
rect 10502 8134 10554 8186
rect 16182 8134 16234 8186
rect 16246 8134 16298 8186
rect 16310 8134 16362 8186
rect 16374 8134 16426 8186
rect 16438 8134 16490 8186
rect 16502 8134 16554 8186
rect 22182 8134 22234 8186
rect 22246 8134 22298 8186
rect 22310 8134 22362 8186
rect 22374 8134 22426 8186
rect 22438 8134 22490 8186
rect 22502 8134 22554 8186
rect 28182 8134 28234 8186
rect 28246 8134 28298 8186
rect 28310 8134 28362 8186
rect 28374 8134 28426 8186
rect 28438 8134 28490 8186
rect 28502 8134 28554 8186
rect 9772 8075 9824 8084
rect 2504 7896 2556 7948
rect 5356 7828 5408 7880
rect 7288 7828 7340 7880
rect 8668 7828 8720 7880
rect 9312 7871 9364 7880
rect 9312 7837 9321 7871
rect 9321 7837 9355 7871
rect 9355 7837 9364 7871
rect 9312 7828 9364 7837
rect 9772 8041 9781 8075
rect 9781 8041 9815 8075
rect 9815 8041 9824 8075
rect 9772 8032 9824 8041
rect 18512 8032 18564 8084
rect 19340 8032 19392 8084
rect 20628 8032 20680 8084
rect 22744 8032 22796 8084
rect 27068 8032 27120 8084
rect 31116 8075 31168 8084
rect 31116 8041 31125 8075
rect 31125 8041 31159 8075
rect 31159 8041 31168 8075
rect 31116 8032 31168 8041
rect 13360 7964 13412 8016
rect 11612 7896 11664 7948
rect 12532 7896 12584 7948
rect 9680 7828 9732 7880
rect 11336 7828 11388 7880
rect 5632 7760 5684 7812
rect 9772 7760 9824 7812
rect 10508 7760 10560 7812
rect 10692 7760 10744 7812
rect 6736 7735 6788 7744
rect 6736 7701 6745 7735
rect 6745 7701 6779 7735
rect 6779 7701 6788 7735
rect 6736 7692 6788 7701
rect 7472 7692 7524 7744
rect 11428 7760 11480 7812
rect 12256 7760 12308 7812
rect 13452 7692 13504 7744
rect 14096 7896 14148 7948
rect 19432 7964 19484 8016
rect 19800 7964 19852 8016
rect 20628 7939 20680 7948
rect 20628 7905 20637 7939
rect 20637 7905 20671 7939
rect 20671 7905 20680 7939
rect 20628 7896 20680 7905
rect 22100 7896 22152 7948
rect 22836 7896 22888 7948
rect 23388 7939 23440 7948
rect 23388 7905 23397 7939
rect 23397 7905 23431 7939
rect 23431 7905 23440 7939
rect 23388 7896 23440 7905
rect 24860 7896 24912 7948
rect 16672 7828 16724 7880
rect 16856 7871 16908 7880
rect 16856 7837 16890 7871
rect 16890 7837 16908 7871
rect 16856 7828 16908 7837
rect 21824 7828 21876 7880
rect 25780 7871 25832 7880
rect 25780 7837 25789 7871
rect 25789 7837 25823 7871
rect 25823 7837 25832 7871
rect 25780 7828 25832 7837
rect 23664 7760 23716 7812
rect 24952 7760 25004 7812
rect 28816 7828 28868 7880
rect 16580 7692 16632 7744
rect 19616 7692 19668 7744
rect 20628 7692 20680 7744
rect 21640 7692 21692 7744
rect 28632 7803 28684 7812
rect 28632 7769 28650 7803
rect 28650 7769 28684 7803
rect 28632 7760 28684 7769
rect 31852 7760 31904 7812
rect 27344 7692 27396 7744
rect 4922 7590 4974 7642
rect 4986 7590 5038 7642
rect 5050 7590 5102 7642
rect 5114 7590 5166 7642
rect 5178 7590 5230 7642
rect 5242 7590 5294 7642
rect 10922 7590 10974 7642
rect 10986 7590 11038 7642
rect 11050 7590 11102 7642
rect 11114 7590 11166 7642
rect 11178 7590 11230 7642
rect 11242 7590 11294 7642
rect 16922 7590 16974 7642
rect 16986 7590 17038 7642
rect 17050 7590 17102 7642
rect 17114 7590 17166 7642
rect 17178 7590 17230 7642
rect 17242 7590 17294 7642
rect 22922 7590 22974 7642
rect 22986 7590 23038 7642
rect 23050 7590 23102 7642
rect 23114 7590 23166 7642
rect 23178 7590 23230 7642
rect 23242 7590 23294 7642
rect 28922 7590 28974 7642
rect 28986 7590 29038 7642
rect 29050 7590 29102 7642
rect 29114 7590 29166 7642
rect 29178 7590 29230 7642
rect 29242 7590 29294 7642
rect 5632 7531 5684 7540
rect 5632 7497 5641 7531
rect 5641 7497 5675 7531
rect 5675 7497 5684 7531
rect 5632 7488 5684 7497
rect 6000 7488 6052 7540
rect 6552 7488 6604 7540
rect 5908 7420 5960 7472
rect 6920 7420 6972 7472
rect 8852 7420 8904 7472
rect 9956 7488 10008 7540
rect 9680 7420 9732 7472
rect 10508 7488 10560 7540
rect 14096 7488 14148 7540
rect 19616 7488 19668 7540
rect 6736 7352 6788 7404
rect 8760 7395 8812 7404
rect 8760 7361 8769 7395
rect 8769 7361 8803 7395
rect 8803 7361 8812 7395
rect 8760 7352 8812 7361
rect 7288 7284 7340 7336
rect 7748 7284 7800 7336
rect 8208 7284 8260 7336
rect 8576 7327 8628 7336
rect 8576 7293 8585 7327
rect 8585 7293 8619 7327
rect 8619 7293 8628 7327
rect 8576 7284 8628 7293
rect 11612 7352 11664 7404
rect 13452 7395 13504 7404
rect 7196 7191 7248 7200
rect 7196 7157 7205 7191
rect 7205 7157 7239 7191
rect 7239 7157 7248 7191
rect 7196 7148 7248 7157
rect 12532 7284 12584 7336
rect 13452 7361 13475 7395
rect 13475 7361 13504 7395
rect 13452 7352 13504 7361
rect 19892 7420 19944 7472
rect 23388 7488 23440 7540
rect 25780 7488 25832 7540
rect 27804 7488 27856 7540
rect 28632 7488 28684 7540
rect 10876 7148 10928 7200
rect 14740 7284 14792 7336
rect 15108 7327 15160 7336
rect 15108 7293 15117 7327
rect 15117 7293 15151 7327
rect 15151 7293 15160 7327
rect 15108 7284 15160 7293
rect 21640 7352 21692 7404
rect 27436 7463 27488 7472
rect 27436 7429 27445 7463
rect 27445 7429 27479 7463
rect 27479 7429 27488 7463
rect 27436 7420 27488 7429
rect 25596 7352 25648 7404
rect 15476 7216 15528 7268
rect 22836 7284 22888 7336
rect 13452 7148 13504 7200
rect 14648 7191 14700 7200
rect 14648 7157 14657 7191
rect 14657 7157 14691 7191
rect 14691 7157 14700 7191
rect 14648 7148 14700 7157
rect 27344 7216 27396 7268
rect 22100 7148 22152 7200
rect 4182 7046 4234 7098
rect 4246 7046 4298 7098
rect 4310 7046 4362 7098
rect 4374 7046 4426 7098
rect 4438 7046 4490 7098
rect 4502 7046 4554 7098
rect 10182 7046 10234 7098
rect 10246 7046 10298 7098
rect 10310 7046 10362 7098
rect 10374 7046 10426 7098
rect 10438 7046 10490 7098
rect 10502 7046 10554 7098
rect 16182 7046 16234 7098
rect 16246 7046 16298 7098
rect 16310 7046 16362 7098
rect 16374 7046 16426 7098
rect 16438 7046 16490 7098
rect 16502 7046 16554 7098
rect 22182 7046 22234 7098
rect 22246 7046 22298 7098
rect 22310 7046 22362 7098
rect 22374 7046 22426 7098
rect 22438 7046 22490 7098
rect 22502 7046 22554 7098
rect 28182 7046 28234 7098
rect 28246 7046 28298 7098
rect 28310 7046 28362 7098
rect 28374 7046 28426 7098
rect 28438 7046 28490 7098
rect 28502 7046 28554 7098
rect 8760 6944 8812 6996
rect 10692 6987 10744 6996
rect 10692 6953 10701 6987
rect 10701 6953 10735 6987
rect 10735 6953 10744 6987
rect 10692 6944 10744 6953
rect 12072 6944 12124 6996
rect 15384 6944 15436 6996
rect 15476 6987 15528 6996
rect 15476 6953 15485 6987
rect 15485 6953 15519 6987
rect 15519 6953 15528 6987
rect 15476 6944 15528 6953
rect 16580 6944 16632 6996
rect 24676 6944 24728 6996
rect 8208 6876 8260 6928
rect 13728 6919 13780 6928
rect 13728 6885 13737 6919
rect 13737 6885 13771 6919
rect 13771 6885 13780 6919
rect 13728 6876 13780 6885
rect 5356 6808 5408 6860
rect 9772 6808 9824 6860
rect 6920 6783 6972 6792
rect 6920 6749 6929 6783
rect 6929 6749 6963 6783
rect 6963 6749 6972 6783
rect 6920 6740 6972 6749
rect 9588 6740 9640 6792
rect 5816 6672 5868 6724
rect 5908 6672 5960 6724
rect 10048 6672 10100 6724
rect 10876 6740 10928 6792
rect 6644 6604 6696 6656
rect 8300 6647 8352 6656
rect 8300 6613 8309 6647
rect 8309 6613 8343 6647
rect 8343 6613 8352 6647
rect 8300 6604 8352 6613
rect 9772 6604 9824 6656
rect 13268 6740 13320 6792
rect 13452 6808 13504 6860
rect 13544 6783 13596 6792
rect 13544 6749 13553 6783
rect 13553 6749 13587 6783
rect 13587 6749 13596 6783
rect 13544 6740 13596 6749
rect 16672 6808 16724 6860
rect 19432 6876 19484 6928
rect 21732 6876 21784 6928
rect 22192 6876 22244 6928
rect 20812 6808 20864 6860
rect 17684 6740 17736 6792
rect 19156 6740 19208 6792
rect 12808 6672 12860 6724
rect 24124 6740 24176 6792
rect 13912 6672 13964 6724
rect 14004 6672 14056 6724
rect 12164 6604 12216 6656
rect 20628 6672 20680 6724
rect 22008 6672 22060 6724
rect 24676 6672 24728 6724
rect 25504 6740 25556 6792
rect 16764 6647 16816 6656
rect 16764 6613 16773 6647
rect 16773 6613 16807 6647
rect 16807 6613 16816 6647
rect 16764 6604 16816 6613
rect 17316 6647 17368 6656
rect 17316 6613 17325 6647
rect 17325 6613 17359 6647
rect 17359 6613 17368 6647
rect 17316 6604 17368 6613
rect 18788 6604 18840 6656
rect 19064 6604 19116 6656
rect 21824 6604 21876 6656
rect 24032 6604 24084 6656
rect 24216 6604 24268 6656
rect 25780 6604 25832 6656
rect 26424 6604 26476 6656
rect 4922 6502 4974 6554
rect 4986 6502 5038 6554
rect 5050 6502 5102 6554
rect 5114 6502 5166 6554
rect 5178 6502 5230 6554
rect 5242 6502 5294 6554
rect 10922 6502 10974 6554
rect 10986 6502 11038 6554
rect 11050 6502 11102 6554
rect 11114 6502 11166 6554
rect 11178 6502 11230 6554
rect 11242 6502 11294 6554
rect 16922 6502 16974 6554
rect 16986 6502 17038 6554
rect 17050 6502 17102 6554
rect 17114 6502 17166 6554
rect 17178 6502 17230 6554
rect 17242 6502 17294 6554
rect 22922 6502 22974 6554
rect 22986 6502 23038 6554
rect 23050 6502 23102 6554
rect 23114 6502 23166 6554
rect 23178 6502 23230 6554
rect 23242 6502 23294 6554
rect 28922 6502 28974 6554
rect 28986 6502 29038 6554
rect 29050 6502 29102 6554
rect 29114 6502 29166 6554
rect 29178 6502 29230 6554
rect 29242 6502 29294 6554
rect 4620 6400 4672 6452
rect 5356 6400 5408 6452
rect 5908 6443 5960 6452
rect 5908 6409 5917 6443
rect 5917 6409 5951 6443
rect 5951 6409 5960 6443
rect 5908 6400 5960 6409
rect 7196 6400 7248 6452
rect 940 6264 992 6316
rect 5448 6264 5500 6316
rect 5724 6307 5776 6316
rect 5724 6273 5733 6307
rect 5733 6273 5767 6307
rect 5767 6273 5776 6307
rect 5724 6264 5776 6273
rect 9220 6400 9272 6452
rect 8300 6264 8352 6316
rect 8576 6307 8628 6316
rect 8576 6273 8585 6307
rect 8585 6273 8619 6307
rect 8619 6273 8628 6307
rect 8576 6264 8628 6273
rect 8484 6196 8536 6248
rect 8852 6307 8904 6316
rect 8852 6273 8861 6307
rect 8861 6273 8895 6307
rect 8895 6273 8904 6307
rect 8852 6264 8904 6273
rect 8944 6307 8996 6316
rect 8944 6273 8953 6307
rect 8953 6273 8987 6307
rect 8987 6273 8996 6307
rect 8944 6264 8996 6273
rect 9588 6264 9640 6316
rect 12256 6400 12308 6452
rect 12532 6400 12584 6452
rect 13268 6332 13320 6384
rect 12164 6264 12216 6316
rect 7472 6128 7524 6180
rect 7840 6103 7892 6112
rect 7840 6069 7849 6103
rect 7849 6069 7883 6103
rect 7883 6069 7892 6103
rect 7840 6060 7892 6069
rect 11704 6103 11756 6112
rect 11704 6069 11713 6103
rect 11713 6069 11747 6103
rect 11747 6069 11756 6103
rect 11704 6060 11756 6069
rect 12072 6060 12124 6112
rect 14004 6443 14056 6452
rect 14004 6409 14013 6443
rect 14013 6409 14047 6443
rect 14047 6409 14056 6443
rect 14004 6400 14056 6409
rect 14648 6400 14700 6452
rect 17684 6443 17736 6452
rect 17684 6409 17693 6443
rect 17693 6409 17727 6443
rect 17727 6409 17736 6443
rect 17684 6400 17736 6409
rect 19156 6400 19208 6452
rect 19524 6443 19576 6452
rect 19524 6409 19533 6443
rect 19533 6409 19567 6443
rect 19567 6409 19576 6443
rect 19524 6400 19576 6409
rect 19708 6400 19760 6452
rect 19064 6332 19116 6384
rect 19248 6375 19300 6384
rect 19248 6341 19253 6375
rect 19253 6341 19287 6375
rect 19287 6341 19300 6375
rect 19248 6332 19300 6341
rect 22008 6375 22060 6384
rect 22008 6341 22017 6375
rect 22017 6341 22051 6375
rect 22051 6341 22060 6375
rect 22008 6332 22060 6341
rect 16764 6196 16816 6248
rect 17868 6239 17920 6248
rect 17868 6205 17877 6239
rect 17877 6205 17911 6239
rect 17911 6205 17920 6239
rect 17868 6196 17920 6205
rect 19386 6307 19438 6316
rect 19386 6273 19395 6307
rect 19395 6273 19429 6307
rect 19429 6273 19438 6307
rect 19386 6264 19438 6273
rect 22100 6307 22152 6316
rect 22100 6273 22109 6307
rect 22109 6273 22143 6307
rect 22143 6273 22152 6307
rect 22100 6264 22152 6273
rect 22192 6307 22244 6316
rect 22192 6273 22201 6307
rect 22201 6273 22235 6307
rect 22235 6273 22244 6307
rect 22192 6264 22244 6273
rect 22652 6400 22704 6452
rect 23756 6400 23808 6452
rect 24124 6400 24176 6452
rect 25596 6375 25648 6384
rect 25596 6341 25605 6375
rect 25605 6341 25639 6375
rect 25639 6341 25648 6375
rect 25596 6332 25648 6341
rect 21548 6239 21600 6248
rect 21548 6205 21557 6239
rect 21557 6205 21591 6239
rect 21591 6205 21600 6239
rect 21548 6196 21600 6205
rect 23664 6239 23716 6248
rect 23664 6205 23673 6239
rect 23673 6205 23707 6239
rect 23707 6205 23716 6239
rect 23664 6196 23716 6205
rect 25504 6128 25556 6180
rect 12808 6060 12860 6112
rect 17408 6060 17460 6112
rect 18236 6060 18288 6112
rect 20996 6103 21048 6112
rect 20996 6069 21005 6103
rect 21005 6069 21039 6103
rect 21039 6069 21048 6103
rect 20996 6060 21048 6069
rect 23572 6060 23624 6112
rect 25780 6060 25832 6112
rect 4182 5958 4234 6010
rect 4246 5958 4298 6010
rect 4310 5958 4362 6010
rect 4374 5958 4426 6010
rect 4438 5958 4490 6010
rect 4502 5958 4554 6010
rect 10182 5958 10234 6010
rect 10246 5958 10298 6010
rect 10310 5958 10362 6010
rect 10374 5958 10426 6010
rect 10438 5958 10490 6010
rect 10502 5958 10554 6010
rect 16182 5958 16234 6010
rect 16246 5958 16298 6010
rect 16310 5958 16362 6010
rect 16374 5958 16426 6010
rect 16438 5958 16490 6010
rect 16502 5958 16554 6010
rect 22182 5958 22234 6010
rect 22246 5958 22298 6010
rect 22310 5958 22362 6010
rect 22374 5958 22426 6010
rect 22438 5958 22490 6010
rect 22502 5958 22554 6010
rect 28182 5958 28234 6010
rect 28246 5958 28298 6010
rect 28310 5958 28362 6010
rect 28374 5958 28426 6010
rect 28438 5958 28490 6010
rect 28502 5958 28554 6010
rect 5724 5856 5776 5908
rect 7840 5856 7892 5908
rect 7748 5720 7800 5772
rect 11612 5856 11664 5908
rect 12808 5899 12860 5908
rect 12808 5865 12817 5899
rect 12817 5865 12851 5899
rect 12851 5865 12860 5899
rect 12808 5856 12860 5865
rect 18236 5899 18288 5908
rect 18236 5865 18245 5899
rect 18245 5865 18279 5899
rect 18279 5865 18288 5899
rect 18236 5856 18288 5865
rect 13912 5720 13964 5772
rect 14280 5720 14332 5772
rect 16672 5720 16724 5772
rect 17868 5720 17920 5772
rect 18788 5763 18840 5772
rect 18788 5729 18797 5763
rect 18797 5729 18831 5763
rect 18831 5729 18840 5763
rect 18788 5720 18840 5729
rect 19248 5720 19300 5772
rect 12164 5652 12216 5704
rect 12808 5652 12860 5704
rect 18880 5652 18932 5704
rect 5356 5584 5408 5636
rect 7472 5584 7524 5636
rect 11704 5627 11756 5636
rect 11704 5593 11738 5627
rect 11738 5593 11756 5627
rect 11704 5584 11756 5593
rect 17316 5584 17368 5636
rect 14096 5559 14148 5568
rect 14096 5525 14105 5559
rect 14105 5525 14139 5559
rect 14139 5525 14148 5559
rect 14096 5516 14148 5525
rect 15108 5516 15160 5568
rect 18328 5559 18380 5568
rect 18328 5525 18337 5559
rect 18337 5525 18371 5559
rect 18371 5525 18380 5559
rect 18328 5516 18380 5525
rect 20996 5856 21048 5908
rect 21824 5856 21876 5908
rect 23572 5856 23624 5908
rect 23756 5856 23808 5908
rect 20628 5763 20680 5772
rect 20628 5729 20637 5763
rect 20637 5729 20671 5763
rect 20671 5729 20680 5763
rect 20628 5720 20680 5729
rect 20812 5763 20864 5772
rect 20812 5729 20821 5763
rect 20821 5729 20855 5763
rect 20855 5729 20864 5763
rect 20812 5720 20864 5729
rect 21640 5720 21692 5772
rect 21916 5763 21968 5772
rect 21916 5729 21925 5763
rect 21925 5729 21959 5763
rect 21959 5729 21968 5763
rect 25780 5831 25832 5840
rect 25780 5797 25789 5831
rect 25789 5797 25823 5831
rect 25823 5797 25832 5831
rect 25780 5788 25832 5797
rect 21916 5720 21968 5729
rect 23664 5720 23716 5772
rect 24032 5652 24084 5704
rect 24216 5652 24268 5704
rect 19708 5516 19760 5568
rect 19800 5516 19852 5568
rect 21272 5559 21324 5568
rect 21272 5525 21281 5559
rect 21281 5525 21315 5559
rect 21315 5525 21324 5559
rect 21272 5516 21324 5525
rect 21640 5559 21692 5568
rect 21640 5525 21649 5559
rect 21649 5525 21683 5559
rect 21683 5525 21692 5559
rect 21640 5516 21692 5525
rect 4922 5414 4974 5466
rect 4986 5414 5038 5466
rect 5050 5414 5102 5466
rect 5114 5414 5166 5466
rect 5178 5414 5230 5466
rect 5242 5414 5294 5466
rect 10922 5414 10974 5466
rect 10986 5414 11038 5466
rect 11050 5414 11102 5466
rect 11114 5414 11166 5466
rect 11178 5414 11230 5466
rect 11242 5414 11294 5466
rect 16922 5414 16974 5466
rect 16986 5414 17038 5466
rect 17050 5414 17102 5466
rect 17114 5414 17166 5466
rect 17178 5414 17230 5466
rect 17242 5414 17294 5466
rect 22922 5414 22974 5466
rect 22986 5414 23038 5466
rect 23050 5414 23102 5466
rect 23114 5414 23166 5466
rect 23178 5414 23230 5466
rect 23242 5414 23294 5466
rect 28922 5414 28974 5466
rect 28986 5414 29038 5466
rect 29050 5414 29102 5466
rect 29114 5414 29166 5466
rect 29178 5414 29230 5466
rect 29242 5414 29294 5466
rect 8668 5312 8720 5364
rect 9772 5312 9824 5364
rect 13912 5312 13964 5364
rect 17316 5312 17368 5364
rect 17408 5312 17460 5364
rect 18880 5355 18932 5364
rect 18880 5321 18889 5355
rect 18889 5321 18923 5355
rect 18923 5321 18932 5355
rect 18880 5312 18932 5321
rect 8024 5219 8076 5228
rect 8024 5185 8033 5219
rect 8033 5185 8067 5219
rect 8067 5185 8076 5219
rect 8024 5176 8076 5185
rect 14280 5244 14332 5296
rect 13084 5219 13136 5228
rect 13084 5185 13118 5219
rect 13118 5185 13136 5219
rect 13084 5176 13136 5185
rect 21272 5312 21324 5364
rect 21640 5312 21692 5364
rect 17776 5219 17828 5228
rect 17776 5185 17810 5219
rect 17810 5185 17828 5219
rect 17776 5176 17828 5185
rect 19800 5176 19852 5228
rect 19892 5219 19944 5228
rect 19892 5185 19901 5219
rect 19901 5185 19935 5219
rect 19935 5185 19944 5219
rect 19892 5176 19944 5185
rect 22100 5176 22152 5228
rect 12808 5151 12860 5160
rect 12808 5117 12817 5151
rect 12817 5117 12851 5151
rect 12851 5117 12860 5151
rect 12808 5108 12860 5117
rect 8852 5040 8904 5092
rect 7288 4972 7340 5024
rect 9220 5015 9272 5024
rect 9220 4981 9229 5015
rect 9229 4981 9263 5015
rect 9263 4981 9272 5015
rect 9220 4972 9272 4981
rect 21548 5040 21600 5092
rect 15476 4972 15528 5024
rect 21364 5015 21416 5024
rect 21364 4981 21373 5015
rect 21373 4981 21407 5015
rect 21407 4981 21416 5015
rect 21364 4972 21416 4981
rect 4182 4870 4234 4922
rect 4246 4870 4298 4922
rect 4310 4870 4362 4922
rect 4374 4870 4426 4922
rect 4438 4870 4490 4922
rect 4502 4870 4554 4922
rect 10182 4870 10234 4922
rect 10246 4870 10298 4922
rect 10310 4870 10362 4922
rect 10374 4870 10426 4922
rect 10438 4870 10490 4922
rect 10502 4870 10554 4922
rect 16182 4870 16234 4922
rect 16246 4870 16298 4922
rect 16310 4870 16362 4922
rect 16374 4870 16426 4922
rect 16438 4870 16490 4922
rect 16502 4870 16554 4922
rect 22182 4870 22234 4922
rect 22246 4870 22298 4922
rect 22310 4870 22362 4922
rect 22374 4870 22426 4922
rect 22438 4870 22490 4922
rect 22502 4870 22554 4922
rect 28182 4870 28234 4922
rect 28246 4870 28298 4922
rect 28310 4870 28362 4922
rect 28374 4870 28426 4922
rect 28438 4870 28490 4922
rect 28502 4870 28554 4922
rect 8024 4768 8076 4820
rect 9220 4768 9272 4820
rect 13084 4768 13136 4820
rect 14096 4768 14148 4820
rect 17776 4768 17828 4820
rect 22100 4811 22152 4820
rect 22100 4777 22109 4811
rect 22109 4777 22143 4811
rect 22143 4777 22152 4811
rect 22100 4768 22152 4777
rect 8852 4700 8904 4752
rect 6920 4632 6972 4684
rect 8392 4632 8444 4684
rect 7288 4564 7340 4616
rect 10784 4564 10836 4616
rect 15200 4632 15252 4684
rect 19892 4632 19944 4684
rect 18328 4564 18380 4616
rect 21364 4564 21416 4616
rect 7288 4471 7340 4480
rect 7288 4437 7297 4471
rect 7297 4437 7331 4471
rect 7331 4437 7340 4471
rect 7288 4428 7340 4437
rect 15476 4496 15528 4548
rect 16580 4496 16632 4548
rect 10508 4471 10560 4480
rect 10508 4437 10517 4471
rect 10517 4437 10551 4471
rect 10551 4437 10560 4471
rect 10508 4428 10560 4437
rect 15016 4428 15068 4480
rect 31208 4428 31260 4480
rect 4922 4326 4974 4378
rect 4986 4326 5038 4378
rect 5050 4326 5102 4378
rect 5114 4326 5166 4378
rect 5178 4326 5230 4378
rect 5242 4326 5294 4378
rect 10922 4326 10974 4378
rect 10986 4326 11038 4378
rect 11050 4326 11102 4378
rect 11114 4326 11166 4378
rect 11178 4326 11230 4378
rect 11242 4326 11294 4378
rect 16922 4326 16974 4378
rect 16986 4326 17038 4378
rect 17050 4326 17102 4378
rect 17114 4326 17166 4378
rect 17178 4326 17230 4378
rect 17242 4326 17294 4378
rect 22922 4326 22974 4378
rect 22986 4326 23038 4378
rect 23050 4326 23102 4378
rect 23114 4326 23166 4378
rect 23178 4326 23230 4378
rect 23242 4326 23294 4378
rect 28922 4326 28974 4378
rect 28986 4326 29038 4378
rect 29050 4326 29102 4378
rect 29114 4326 29166 4378
rect 29178 4326 29230 4378
rect 29242 4326 29294 4378
rect 7288 4224 7340 4276
rect 8392 4224 8444 4276
rect 10508 4224 10560 4276
rect 15016 4267 15068 4276
rect 15016 4233 15025 4267
rect 15025 4233 15059 4267
rect 15059 4233 15068 4267
rect 15016 4224 15068 4233
rect 17408 4156 17460 4208
rect 6920 4088 6972 4140
rect 10048 4020 10100 4072
rect 10600 4088 10652 4140
rect 15292 4088 15344 4140
rect 15660 4088 15712 4140
rect 10692 4020 10744 4072
rect 11888 4020 11940 4072
rect 14648 3952 14700 4004
rect 9680 3927 9732 3936
rect 9680 3893 9689 3927
rect 9689 3893 9723 3927
rect 9723 3893 9732 3927
rect 9680 3884 9732 3893
rect 10048 3884 10100 3936
rect 15384 3927 15436 3936
rect 15384 3893 15393 3927
rect 15393 3893 15427 3927
rect 15427 3893 15436 3927
rect 15384 3884 15436 3893
rect 15568 3884 15620 3936
rect 4182 3782 4234 3834
rect 4246 3782 4298 3834
rect 4310 3782 4362 3834
rect 4374 3782 4426 3834
rect 4438 3782 4490 3834
rect 4502 3782 4554 3834
rect 10182 3782 10234 3834
rect 10246 3782 10298 3834
rect 10310 3782 10362 3834
rect 10374 3782 10426 3834
rect 10438 3782 10490 3834
rect 10502 3782 10554 3834
rect 16182 3782 16234 3834
rect 16246 3782 16298 3834
rect 16310 3782 16362 3834
rect 16374 3782 16426 3834
rect 16438 3782 16490 3834
rect 16502 3782 16554 3834
rect 22182 3782 22234 3834
rect 22246 3782 22298 3834
rect 22310 3782 22362 3834
rect 22374 3782 22426 3834
rect 22438 3782 22490 3834
rect 22502 3782 22554 3834
rect 28182 3782 28234 3834
rect 28246 3782 28298 3834
rect 28310 3782 28362 3834
rect 28374 3782 28426 3834
rect 28438 3782 28490 3834
rect 28502 3782 28554 3834
rect 9680 3680 9732 3732
rect 10048 3680 10100 3732
rect 9772 3476 9824 3528
rect 12164 3587 12216 3596
rect 12164 3553 12173 3587
rect 12173 3553 12207 3587
rect 12207 3553 12216 3587
rect 12164 3544 12216 3553
rect 14556 3587 14608 3596
rect 14556 3553 14565 3587
rect 14565 3553 14599 3587
rect 14599 3553 14608 3587
rect 14556 3544 14608 3553
rect 14648 3587 14700 3596
rect 14648 3553 14657 3587
rect 14657 3553 14691 3587
rect 14691 3553 14700 3587
rect 14648 3544 14700 3553
rect 15384 3680 15436 3732
rect 15568 3680 15620 3732
rect 17408 3723 17460 3732
rect 17408 3689 17417 3723
rect 17417 3689 17451 3723
rect 17451 3689 17460 3723
rect 17408 3680 17460 3689
rect 17868 3680 17920 3732
rect 15200 3612 15252 3664
rect 15476 3544 15528 3596
rect 9036 3408 9088 3460
rect 9496 3383 9548 3392
rect 9496 3349 9505 3383
rect 9505 3349 9539 3383
rect 9539 3349 9548 3383
rect 9496 3340 9548 3349
rect 9864 3383 9916 3392
rect 9864 3349 9873 3383
rect 9873 3349 9907 3383
rect 9907 3349 9916 3383
rect 9864 3340 9916 3349
rect 11612 3408 11664 3460
rect 12440 3451 12492 3460
rect 12440 3417 12449 3451
rect 12449 3417 12483 3451
rect 12483 3417 12492 3451
rect 12440 3408 12492 3417
rect 13728 3408 13780 3460
rect 11888 3340 11940 3392
rect 13912 3383 13964 3392
rect 13912 3349 13921 3383
rect 13921 3349 13955 3383
rect 13955 3349 13964 3383
rect 13912 3340 13964 3349
rect 14096 3383 14148 3392
rect 14096 3349 14105 3383
rect 14105 3349 14139 3383
rect 14139 3349 14148 3383
rect 14096 3340 14148 3349
rect 16672 3408 16724 3460
rect 4922 3238 4974 3290
rect 4986 3238 5038 3290
rect 5050 3238 5102 3290
rect 5114 3238 5166 3290
rect 5178 3238 5230 3290
rect 5242 3238 5294 3290
rect 10922 3238 10974 3290
rect 10986 3238 11038 3290
rect 11050 3238 11102 3290
rect 11114 3238 11166 3290
rect 11178 3238 11230 3290
rect 11242 3238 11294 3290
rect 16922 3238 16974 3290
rect 16986 3238 17038 3290
rect 17050 3238 17102 3290
rect 17114 3238 17166 3290
rect 17178 3238 17230 3290
rect 17242 3238 17294 3290
rect 22922 3238 22974 3290
rect 22986 3238 23038 3290
rect 23050 3238 23102 3290
rect 23114 3238 23166 3290
rect 23178 3238 23230 3290
rect 23242 3238 23294 3290
rect 28922 3238 28974 3290
rect 28986 3238 29038 3290
rect 29050 3238 29102 3290
rect 29114 3238 29166 3290
rect 29178 3238 29230 3290
rect 29242 3238 29294 3290
rect 9496 3136 9548 3188
rect 10784 3179 10836 3188
rect 10784 3145 10793 3179
rect 10793 3145 10827 3179
rect 10827 3145 10836 3179
rect 10784 3136 10836 3145
rect 11612 3179 11664 3188
rect 11612 3145 11621 3179
rect 11621 3145 11655 3179
rect 11655 3145 11664 3179
rect 11612 3136 11664 3145
rect 12440 3136 12492 3188
rect 13728 3179 13780 3188
rect 13728 3145 13737 3179
rect 13737 3145 13771 3179
rect 13771 3145 13780 3179
rect 13728 3136 13780 3145
rect 14096 3136 14148 3188
rect 16580 3136 16632 3188
rect 16672 3136 16724 3188
rect 9864 3068 9916 3120
rect 6920 3000 6972 3052
rect 9036 3043 9088 3052
rect 9036 3009 9045 3043
rect 9045 3009 9079 3043
rect 9079 3009 9088 3043
rect 9036 3000 9088 3009
rect 9772 2932 9824 2984
rect 4182 2694 4234 2746
rect 4246 2694 4298 2746
rect 4310 2694 4362 2746
rect 4374 2694 4426 2746
rect 4438 2694 4490 2746
rect 4502 2694 4554 2746
rect 10182 2694 10234 2746
rect 10246 2694 10298 2746
rect 10310 2694 10362 2746
rect 10374 2694 10426 2746
rect 10438 2694 10490 2746
rect 10502 2694 10554 2746
rect 16182 2694 16234 2746
rect 16246 2694 16298 2746
rect 16310 2694 16362 2746
rect 16374 2694 16426 2746
rect 16438 2694 16490 2746
rect 16502 2694 16554 2746
rect 22182 2694 22234 2746
rect 22246 2694 22298 2746
rect 22310 2694 22362 2746
rect 22374 2694 22426 2746
rect 22438 2694 22490 2746
rect 22502 2694 22554 2746
rect 28182 2694 28234 2746
rect 28246 2694 28298 2746
rect 28310 2694 28362 2746
rect 28374 2694 28426 2746
rect 28438 2694 28490 2746
rect 28502 2694 28554 2746
rect 29368 2592 29420 2644
rect 13912 2456 13964 2508
rect 11888 2431 11940 2440
rect 11888 2397 11897 2431
rect 11897 2397 11931 2431
rect 11931 2397 11940 2431
rect 11888 2388 11940 2397
rect 17040 2388 17092 2440
rect 17868 2388 17920 2440
rect 29368 2388 29420 2440
rect 31208 2431 31260 2440
rect 31208 2397 31217 2431
rect 31217 2397 31251 2431
rect 31251 2397 31260 2431
rect 31208 2388 31260 2397
rect 20 2320 72 2372
rect 10784 2320 10836 2372
rect 5816 2295 5868 2304
rect 5816 2261 5825 2295
rect 5825 2261 5859 2295
rect 5859 2261 5868 2295
rect 5816 2252 5868 2261
rect 11612 2295 11664 2304
rect 11612 2261 11621 2295
rect 11621 2261 11655 2295
rect 11655 2261 11664 2295
rect 11612 2252 11664 2261
rect 17408 2252 17460 2304
rect 23480 2295 23532 2304
rect 23480 2261 23489 2295
rect 23489 2261 23523 2295
rect 23523 2261 23532 2295
rect 23480 2252 23532 2261
rect 31392 2295 31444 2304
rect 31392 2261 31401 2295
rect 31401 2261 31435 2295
rect 31435 2261 31444 2295
rect 31392 2252 31444 2261
rect 4922 2150 4974 2202
rect 4986 2150 5038 2202
rect 5050 2150 5102 2202
rect 5114 2150 5166 2202
rect 5178 2150 5230 2202
rect 5242 2150 5294 2202
rect 10922 2150 10974 2202
rect 10986 2150 11038 2202
rect 11050 2150 11102 2202
rect 11114 2150 11166 2202
rect 11178 2150 11230 2202
rect 11242 2150 11294 2202
rect 16922 2150 16974 2202
rect 16986 2150 17038 2202
rect 17050 2150 17102 2202
rect 17114 2150 17166 2202
rect 17178 2150 17230 2202
rect 17242 2150 17294 2202
rect 22922 2150 22974 2202
rect 22986 2150 23038 2202
rect 23050 2150 23102 2202
rect 23114 2150 23166 2202
rect 23178 2150 23230 2202
rect 23242 2150 23294 2202
rect 28922 2150 28974 2202
rect 28986 2150 29038 2202
rect 29050 2150 29102 2202
rect 29114 2150 29166 2202
rect 29178 2150 29230 2202
rect 29242 2150 29294 2202
<< metal2 >>
rect 1306 34318 1362 35118
rect 7102 34318 7158 35118
rect 12898 34318 12954 35118
rect 18694 34318 18750 35118
rect 24490 34318 24546 35118
rect 30286 34318 30342 35118
rect 1320 32570 1348 34318
rect 4920 32668 5296 32677
rect 4976 32666 5000 32668
rect 5056 32666 5080 32668
rect 5136 32666 5160 32668
rect 5216 32666 5240 32668
rect 4976 32614 4986 32666
rect 5230 32614 5240 32666
rect 4976 32612 5000 32614
rect 5056 32612 5080 32614
rect 5136 32612 5160 32614
rect 5216 32612 5240 32614
rect 4920 32603 5296 32612
rect 1308 32564 1360 32570
rect 1308 32506 1360 32512
rect 7116 32434 7144 34318
rect 10920 32668 11296 32677
rect 10976 32666 11000 32668
rect 11056 32666 11080 32668
rect 11136 32666 11160 32668
rect 11216 32666 11240 32668
rect 10976 32614 10986 32666
rect 11230 32614 11240 32666
rect 10976 32612 11000 32614
rect 11056 32612 11080 32614
rect 11136 32612 11160 32614
rect 11216 32612 11240 32614
rect 10920 32603 11296 32612
rect 12912 32434 12940 34318
rect 16920 32668 17296 32677
rect 16976 32666 17000 32668
rect 17056 32666 17080 32668
rect 17136 32666 17160 32668
rect 17216 32666 17240 32668
rect 16976 32614 16986 32666
rect 17230 32614 17240 32666
rect 16976 32612 17000 32614
rect 17056 32612 17080 32614
rect 17136 32612 17160 32614
rect 17216 32612 17240 32614
rect 16920 32603 17296 32612
rect 18708 32570 18736 34318
rect 22920 32668 23296 32677
rect 22976 32666 23000 32668
rect 23056 32666 23080 32668
rect 23136 32666 23160 32668
rect 23216 32666 23240 32668
rect 22976 32614 22986 32666
rect 23230 32614 23240 32666
rect 22976 32612 23000 32614
rect 23056 32612 23080 32614
rect 23136 32612 23160 32614
rect 23216 32612 23240 32614
rect 22920 32603 23296 32612
rect 24504 32570 24532 34318
rect 28920 32668 29296 32677
rect 28976 32666 29000 32668
rect 29056 32666 29080 32668
rect 29136 32666 29160 32668
rect 29216 32666 29240 32668
rect 28976 32614 28986 32666
rect 29230 32614 29240 32666
rect 28976 32612 29000 32614
rect 29056 32612 29080 32614
rect 29136 32612 29160 32614
rect 29216 32612 29240 32614
rect 28920 32603 29296 32612
rect 18696 32564 18748 32570
rect 18696 32506 18748 32512
rect 24492 32564 24544 32570
rect 24492 32506 24544 32512
rect 30300 32434 30328 34318
rect 7104 32428 7156 32434
rect 7104 32370 7156 32376
rect 12900 32428 12952 32434
rect 12900 32370 12952 32376
rect 19340 32428 19392 32434
rect 19340 32370 19392 32376
rect 24676 32428 24728 32434
rect 24676 32370 24728 32376
rect 30288 32428 30340 32434
rect 30288 32370 30340 32376
rect 12440 32292 12492 32298
rect 12440 32234 12492 32240
rect 7380 32224 7432 32230
rect 7380 32166 7432 32172
rect 4180 32124 4556 32133
rect 4236 32122 4260 32124
rect 4316 32122 4340 32124
rect 4396 32122 4420 32124
rect 4476 32122 4500 32124
rect 4236 32070 4246 32122
rect 4490 32070 4500 32122
rect 4236 32068 4260 32070
rect 4316 32068 4340 32070
rect 4396 32068 4420 32070
rect 4476 32068 4500 32070
rect 4180 32059 4556 32068
rect 4920 31580 5296 31589
rect 4976 31578 5000 31580
rect 5056 31578 5080 31580
rect 5136 31578 5160 31580
rect 5216 31578 5240 31580
rect 4976 31526 4986 31578
rect 5230 31526 5240 31578
rect 4976 31524 5000 31526
rect 5056 31524 5080 31526
rect 5136 31524 5160 31526
rect 5216 31524 5240 31526
rect 4920 31515 5296 31524
rect 4180 31036 4556 31045
rect 4236 31034 4260 31036
rect 4316 31034 4340 31036
rect 4396 31034 4420 31036
rect 4476 31034 4500 31036
rect 4236 30982 4246 31034
rect 4490 30982 4500 31034
rect 4236 30980 4260 30982
rect 4316 30980 4340 30982
rect 4396 30980 4420 30982
rect 4476 30980 4500 30982
rect 4180 30971 4556 30980
rect 940 30728 992 30734
rect 938 30696 940 30705
rect 992 30696 994 30705
rect 938 30631 994 30640
rect 1584 30592 1636 30598
rect 1584 30534 1636 30540
rect 1596 26234 1624 30534
rect 4920 30492 5296 30501
rect 4976 30490 5000 30492
rect 5056 30490 5080 30492
rect 5136 30490 5160 30492
rect 5216 30490 5240 30492
rect 4976 30438 4986 30490
rect 5230 30438 5240 30490
rect 4976 30436 5000 30438
rect 5056 30436 5080 30438
rect 5136 30436 5160 30438
rect 5216 30436 5240 30438
rect 4920 30427 5296 30436
rect 4180 29948 4556 29957
rect 4236 29946 4260 29948
rect 4316 29946 4340 29948
rect 4396 29946 4420 29948
rect 4476 29946 4500 29948
rect 4236 29894 4246 29946
rect 4490 29894 4500 29946
rect 4236 29892 4260 29894
rect 4316 29892 4340 29894
rect 4396 29892 4420 29894
rect 4476 29892 4500 29894
rect 4180 29883 4556 29892
rect 4920 29404 5296 29413
rect 4976 29402 5000 29404
rect 5056 29402 5080 29404
rect 5136 29402 5160 29404
rect 5216 29402 5240 29404
rect 4976 29350 4986 29402
rect 5230 29350 5240 29402
rect 4976 29348 5000 29350
rect 5056 29348 5080 29350
rect 5136 29348 5160 29350
rect 5216 29348 5240 29350
rect 4920 29339 5296 29348
rect 4180 28860 4556 28869
rect 4236 28858 4260 28860
rect 4316 28858 4340 28860
rect 4396 28858 4420 28860
rect 4476 28858 4500 28860
rect 4236 28806 4246 28858
rect 4490 28806 4500 28858
rect 4236 28804 4260 28806
rect 4316 28804 4340 28806
rect 4396 28804 4420 28806
rect 4476 28804 4500 28806
rect 4180 28795 4556 28804
rect 4920 28316 5296 28325
rect 4976 28314 5000 28316
rect 5056 28314 5080 28316
rect 5136 28314 5160 28316
rect 5216 28314 5240 28316
rect 4976 28262 4986 28314
rect 5230 28262 5240 28314
rect 4976 28260 5000 28262
rect 5056 28260 5080 28262
rect 5136 28260 5160 28262
rect 5216 28260 5240 28262
rect 4920 28251 5296 28260
rect 4180 27772 4556 27781
rect 4236 27770 4260 27772
rect 4316 27770 4340 27772
rect 4396 27770 4420 27772
rect 4476 27770 4500 27772
rect 4236 27718 4246 27770
rect 4490 27718 4500 27770
rect 4236 27716 4260 27718
rect 4316 27716 4340 27718
rect 4396 27716 4420 27718
rect 4476 27716 4500 27718
rect 4180 27707 4556 27716
rect 4804 27396 4856 27402
rect 4804 27338 4856 27344
rect 4180 26684 4556 26693
rect 4236 26682 4260 26684
rect 4316 26682 4340 26684
rect 4396 26682 4420 26684
rect 4476 26682 4500 26684
rect 4236 26630 4246 26682
rect 4490 26630 4500 26682
rect 4236 26628 4260 26630
rect 4316 26628 4340 26630
rect 4396 26628 4420 26630
rect 4476 26628 4500 26630
rect 4180 26619 4556 26628
rect 3976 26240 4028 26246
rect 1596 26206 1716 26234
rect 940 24744 992 24750
rect 940 24686 992 24692
rect 952 24585 980 24686
rect 938 24576 994 24585
rect 938 24511 994 24520
rect 940 18760 992 18766
rect 940 18702 992 18708
rect 952 18465 980 18702
rect 938 18456 994 18465
rect 938 18391 994 18400
rect 1688 14958 1716 26206
rect 3976 26182 4028 26188
rect 3988 25362 4016 26182
rect 4816 25838 4844 27338
rect 4920 27228 5296 27237
rect 4976 27226 5000 27228
rect 5056 27226 5080 27228
rect 5136 27226 5160 27228
rect 5216 27226 5240 27228
rect 4976 27174 4986 27226
rect 5230 27174 5240 27226
rect 4976 27172 5000 27174
rect 5056 27172 5080 27174
rect 5136 27172 5160 27174
rect 5216 27172 5240 27174
rect 4920 27163 5296 27172
rect 6092 26988 6144 26994
rect 6092 26930 6144 26936
rect 4920 26140 5296 26149
rect 4976 26138 5000 26140
rect 5056 26138 5080 26140
rect 5136 26138 5160 26140
rect 5216 26138 5240 26140
rect 4976 26086 4986 26138
rect 5230 26086 5240 26138
rect 4976 26084 5000 26086
rect 5056 26084 5080 26086
rect 5136 26084 5160 26086
rect 5216 26084 5240 26086
rect 4920 26075 5296 26084
rect 5908 25968 5960 25974
rect 5908 25910 5960 25916
rect 4804 25832 4856 25838
rect 4804 25774 4856 25780
rect 4620 25696 4672 25702
rect 4620 25638 4672 25644
rect 4180 25596 4556 25605
rect 4236 25594 4260 25596
rect 4316 25594 4340 25596
rect 4396 25594 4420 25596
rect 4476 25594 4500 25596
rect 4236 25542 4246 25594
rect 4490 25542 4500 25594
rect 4236 25540 4260 25542
rect 4316 25540 4340 25542
rect 4396 25540 4420 25542
rect 4476 25540 4500 25542
rect 4180 25531 4556 25540
rect 3976 25356 4028 25362
rect 3976 25298 4028 25304
rect 3988 24818 4016 25298
rect 4632 24886 4660 25638
rect 4816 25378 4844 25774
rect 5448 25764 5500 25770
rect 5448 25706 5500 25712
rect 5460 25498 5488 25706
rect 5540 25696 5592 25702
rect 5540 25638 5592 25644
rect 5448 25492 5500 25498
rect 5448 25434 5500 25440
rect 4724 25350 4844 25378
rect 4620 24880 4672 24886
rect 4620 24822 4672 24828
rect 3976 24812 4028 24818
rect 3976 24754 4028 24760
rect 3792 24744 3844 24750
rect 3792 24686 3844 24692
rect 3804 23866 3832 24686
rect 4180 24508 4556 24517
rect 4236 24506 4260 24508
rect 4316 24506 4340 24508
rect 4396 24506 4420 24508
rect 4476 24506 4500 24508
rect 4236 24454 4246 24506
rect 4490 24454 4500 24506
rect 4236 24452 4260 24454
rect 4316 24452 4340 24454
rect 4396 24452 4420 24454
rect 4476 24452 4500 24454
rect 4180 24443 4556 24452
rect 3792 23860 3844 23866
rect 3792 23802 3844 23808
rect 4180 23420 4556 23429
rect 4236 23418 4260 23420
rect 4316 23418 4340 23420
rect 4396 23418 4420 23420
rect 4476 23418 4500 23420
rect 4236 23366 4246 23418
rect 4490 23366 4500 23418
rect 4236 23364 4260 23366
rect 4316 23364 4340 23366
rect 4396 23364 4420 23366
rect 4476 23364 4500 23366
rect 4180 23355 4556 23364
rect 4724 23202 4752 25350
rect 4804 25220 4856 25226
rect 4804 25162 4856 25168
rect 4816 24954 4844 25162
rect 4920 25052 5296 25061
rect 4976 25050 5000 25052
rect 5056 25050 5080 25052
rect 5136 25050 5160 25052
rect 5216 25050 5240 25052
rect 4976 24998 4986 25050
rect 5230 24998 5240 25050
rect 4976 24996 5000 24998
rect 5056 24996 5080 24998
rect 5136 24996 5160 24998
rect 5216 24996 5240 24998
rect 4920 24987 5296 24996
rect 5552 24954 5580 25638
rect 5632 25424 5684 25430
rect 5632 25366 5684 25372
rect 4804 24948 4856 24954
rect 4804 24890 4856 24896
rect 5540 24948 5592 24954
rect 5540 24890 5592 24896
rect 5644 24206 5672 25366
rect 5920 25362 5948 25910
rect 6000 25832 6052 25838
rect 6000 25774 6052 25780
rect 6012 25498 6040 25774
rect 6000 25492 6052 25498
rect 6000 25434 6052 25440
rect 6104 25378 6132 26930
rect 6736 26784 6788 26790
rect 6736 26726 6788 26732
rect 6748 26042 6776 26726
rect 7288 26376 7340 26382
rect 7288 26318 7340 26324
rect 7104 26308 7156 26314
rect 7104 26250 7156 26256
rect 7116 26042 7144 26250
rect 6736 26036 6788 26042
rect 6736 25978 6788 25984
rect 7104 26036 7156 26042
rect 7104 25978 7156 25984
rect 6012 25362 6132 25378
rect 5908 25356 5960 25362
rect 5908 25298 5960 25304
rect 6000 25356 6132 25362
rect 6052 25350 6132 25356
rect 6000 25298 6052 25304
rect 5632 24200 5684 24206
rect 5632 24142 5684 24148
rect 5908 24200 5960 24206
rect 5908 24142 5960 24148
rect 5724 24132 5776 24138
rect 5724 24074 5776 24080
rect 4920 23964 5296 23973
rect 4976 23962 5000 23964
rect 5056 23962 5080 23964
rect 5136 23962 5160 23964
rect 5216 23962 5240 23964
rect 4976 23910 4986 23962
rect 5230 23910 5240 23962
rect 4976 23908 5000 23910
rect 5056 23908 5080 23910
rect 5136 23908 5160 23910
rect 5216 23908 5240 23910
rect 4920 23899 5296 23908
rect 4632 23174 4752 23202
rect 4068 22976 4120 22982
rect 4068 22918 4120 22924
rect 3608 22568 3660 22574
rect 3608 22510 3660 22516
rect 3620 22030 3648 22510
rect 3608 22024 3660 22030
rect 3608 21966 3660 21972
rect 4080 21962 4108 22918
rect 4632 22574 4660 23174
rect 4712 23112 4764 23118
rect 4712 23054 4764 23060
rect 4620 22568 4672 22574
rect 4620 22510 4672 22516
rect 4180 22332 4556 22341
rect 4236 22330 4260 22332
rect 4316 22330 4340 22332
rect 4396 22330 4420 22332
rect 4476 22330 4500 22332
rect 4236 22278 4246 22330
rect 4490 22278 4500 22330
rect 4236 22276 4260 22278
rect 4316 22276 4340 22278
rect 4396 22276 4420 22278
rect 4476 22276 4500 22278
rect 4180 22267 4556 22276
rect 4068 21956 4120 21962
rect 4068 21898 4120 21904
rect 4180 21244 4556 21253
rect 4236 21242 4260 21244
rect 4316 21242 4340 21244
rect 4396 21242 4420 21244
rect 4476 21242 4500 21244
rect 4236 21190 4246 21242
rect 4490 21190 4500 21242
rect 4236 21188 4260 21190
rect 4316 21188 4340 21190
rect 4396 21188 4420 21190
rect 4476 21188 4500 21190
rect 4180 21179 4556 21188
rect 4180 20156 4556 20165
rect 4236 20154 4260 20156
rect 4316 20154 4340 20156
rect 4396 20154 4420 20156
rect 4476 20154 4500 20156
rect 4236 20102 4246 20154
rect 4490 20102 4500 20154
rect 4236 20100 4260 20102
rect 4316 20100 4340 20102
rect 4396 20100 4420 20102
rect 4476 20100 4500 20102
rect 4180 20091 4556 20100
rect 3148 19712 3200 19718
rect 3148 19654 3200 19660
rect 3056 19372 3108 19378
rect 3056 19314 3108 19320
rect 3068 18970 3096 19314
rect 3056 18964 3108 18970
rect 3056 18906 3108 18912
rect 3160 18766 3188 19654
rect 3976 19372 4028 19378
rect 3976 19314 4028 19320
rect 4252 19372 4304 19378
rect 4252 19314 4304 19320
rect 3148 18760 3200 18766
rect 3148 18702 3200 18708
rect 3700 18624 3752 18630
rect 3700 18566 3752 18572
rect 3516 17196 3568 17202
rect 3516 17138 3568 17144
rect 3528 16794 3556 17138
rect 3516 16788 3568 16794
rect 3516 16730 3568 16736
rect 3424 16584 3476 16590
rect 3424 16526 3476 16532
rect 3436 16250 3464 16526
rect 3424 16244 3476 16250
rect 3424 16186 3476 16192
rect 1676 14952 1728 14958
rect 1676 14894 1728 14900
rect 2688 14816 2740 14822
rect 2688 14758 2740 14764
rect 3516 14816 3568 14822
rect 3516 14758 3568 14764
rect 2320 14272 2372 14278
rect 2320 14214 2372 14220
rect 2332 13938 2360 14214
rect 2700 14074 2728 14758
rect 3528 14346 3556 14758
rect 3240 14340 3292 14346
rect 3240 14282 3292 14288
rect 3516 14340 3568 14346
rect 3516 14282 3568 14288
rect 2688 14068 2740 14074
rect 2688 14010 2740 14016
rect 2320 13932 2372 13938
rect 2320 13874 2372 13880
rect 3252 13530 3280 14282
rect 3608 14272 3660 14278
rect 3608 14214 3660 14220
rect 3620 14074 3648 14214
rect 3608 14068 3660 14074
rect 3608 14010 3660 14016
rect 3240 13524 3292 13530
rect 3240 13466 3292 13472
rect 1492 12640 1544 12646
rect 1492 12582 1544 12588
rect 1504 12345 1532 12582
rect 1490 12336 1546 12345
rect 1490 12271 1546 12280
rect 2596 11756 2648 11762
rect 2596 11698 2648 11704
rect 2608 11354 2636 11698
rect 3712 11694 3740 18566
rect 3988 17202 4016 19314
rect 4264 19258 4292 19314
rect 4080 19230 4292 19258
rect 4080 18970 4108 19230
rect 4180 19068 4556 19077
rect 4236 19066 4260 19068
rect 4316 19066 4340 19068
rect 4396 19066 4420 19068
rect 4476 19066 4500 19068
rect 4236 19014 4246 19066
rect 4490 19014 4500 19066
rect 4236 19012 4260 19014
rect 4316 19012 4340 19014
rect 4396 19012 4420 19014
rect 4476 19012 4500 19014
rect 4180 19003 4556 19012
rect 4068 18964 4120 18970
rect 4068 18906 4120 18912
rect 4632 18834 4660 22510
rect 4724 22234 4752 23054
rect 5736 23050 5764 24074
rect 5724 23044 5776 23050
rect 5724 22986 5776 22992
rect 4804 22976 4856 22982
rect 4804 22918 4856 22924
rect 5448 22976 5500 22982
rect 5448 22918 5500 22924
rect 4816 22778 4844 22918
rect 4920 22876 5296 22885
rect 4976 22874 5000 22876
rect 5056 22874 5080 22876
rect 5136 22874 5160 22876
rect 5216 22874 5240 22876
rect 4976 22822 4986 22874
rect 5230 22822 5240 22874
rect 4976 22820 5000 22822
rect 5056 22820 5080 22822
rect 5136 22820 5160 22822
rect 5216 22820 5240 22822
rect 4920 22811 5296 22820
rect 5460 22778 5488 22918
rect 4804 22772 4856 22778
rect 4804 22714 4856 22720
rect 5448 22772 5500 22778
rect 5448 22714 5500 22720
rect 5356 22704 5408 22710
rect 5356 22646 5408 22652
rect 4712 22228 4764 22234
rect 4712 22170 4764 22176
rect 5368 22030 5396 22646
rect 5540 22568 5592 22574
rect 5540 22510 5592 22516
rect 5356 22024 5408 22030
rect 5356 21966 5408 21972
rect 4920 21788 5296 21797
rect 4976 21786 5000 21788
rect 5056 21786 5080 21788
rect 5136 21786 5160 21788
rect 5216 21786 5240 21788
rect 4976 21734 4986 21786
rect 5230 21734 5240 21786
rect 4976 21732 5000 21734
rect 5056 21732 5080 21734
rect 5136 21732 5160 21734
rect 5216 21732 5240 21734
rect 4920 21723 5296 21732
rect 5368 21690 5396 21966
rect 5356 21684 5408 21690
rect 5356 21626 5408 21632
rect 5552 21622 5580 22510
rect 5632 21888 5684 21894
rect 5632 21830 5684 21836
rect 5540 21616 5592 21622
rect 5540 21558 5592 21564
rect 5644 21146 5672 21830
rect 5632 21140 5684 21146
rect 5632 21082 5684 21088
rect 4920 20700 5296 20709
rect 4976 20698 5000 20700
rect 5056 20698 5080 20700
rect 5136 20698 5160 20700
rect 5216 20698 5240 20700
rect 4976 20646 4986 20698
rect 5230 20646 5240 20698
rect 4976 20644 5000 20646
rect 5056 20644 5080 20646
rect 5136 20644 5160 20646
rect 5216 20644 5240 20646
rect 4920 20635 5296 20644
rect 4712 19916 4764 19922
rect 4712 19858 4764 19864
rect 4620 18828 4672 18834
rect 4620 18770 4672 18776
rect 4180 17980 4556 17989
rect 4236 17978 4260 17980
rect 4316 17978 4340 17980
rect 4396 17978 4420 17980
rect 4476 17978 4500 17980
rect 4236 17926 4246 17978
rect 4490 17926 4500 17978
rect 4236 17924 4260 17926
rect 4316 17924 4340 17926
rect 4396 17924 4420 17926
rect 4476 17924 4500 17926
rect 4180 17915 4556 17924
rect 3976 17196 4028 17202
rect 3976 17138 4028 17144
rect 3988 16794 4016 17138
rect 4632 17134 4660 18770
rect 4620 17128 4672 17134
rect 4620 17070 4672 17076
rect 4180 16892 4556 16901
rect 4236 16890 4260 16892
rect 4316 16890 4340 16892
rect 4396 16890 4420 16892
rect 4476 16890 4500 16892
rect 4236 16838 4246 16890
rect 4490 16838 4500 16890
rect 4236 16836 4260 16838
rect 4316 16836 4340 16838
rect 4396 16836 4420 16838
rect 4476 16836 4500 16838
rect 4180 16827 4556 16836
rect 3976 16788 4028 16794
rect 3976 16730 4028 16736
rect 4632 16674 4660 17070
rect 4724 16776 4752 19858
rect 5540 19848 5592 19854
rect 5540 19790 5592 19796
rect 4896 19712 4948 19718
rect 4816 19672 4896 19700
rect 4816 18630 4844 19672
rect 4896 19654 4948 19660
rect 4920 19612 5296 19621
rect 4976 19610 5000 19612
rect 5056 19610 5080 19612
rect 5136 19610 5160 19612
rect 5216 19610 5240 19612
rect 4976 19558 4986 19610
rect 5230 19558 5240 19610
rect 4976 19556 5000 19558
rect 5056 19556 5080 19558
rect 5136 19556 5160 19558
rect 5216 19556 5240 19558
rect 4920 19547 5296 19556
rect 5552 19514 5580 19790
rect 5172 19508 5224 19514
rect 5172 19450 5224 19456
rect 5540 19508 5592 19514
rect 5540 19450 5592 19456
rect 5184 18834 5212 19450
rect 5552 18970 5580 19450
rect 5540 18964 5592 18970
rect 5540 18906 5592 18912
rect 5172 18828 5224 18834
rect 5172 18770 5224 18776
rect 5736 18714 5764 22986
rect 5920 22982 5948 24142
rect 5908 22976 5960 22982
rect 5908 22918 5960 22924
rect 5816 22160 5868 22166
rect 5816 22102 5868 22108
rect 5828 19922 5856 22102
rect 5816 19916 5868 19922
rect 5816 19858 5868 19864
rect 5920 19258 5948 22918
rect 6012 22166 6040 25298
rect 7300 25294 7328 26318
rect 6920 25288 6972 25294
rect 6920 25230 6972 25236
rect 7288 25288 7340 25294
rect 7288 25230 7340 25236
rect 6932 24682 6960 25230
rect 6920 24676 6972 24682
rect 6920 24618 6972 24624
rect 6932 24138 6960 24618
rect 6920 24132 6972 24138
rect 6920 24074 6972 24080
rect 6276 23044 6328 23050
rect 6276 22986 6328 22992
rect 6000 22160 6052 22166
rect 6000 22102 6052 22108
rect 6288 21894 6316 22986
rect 7288 22636 7340 22642
rect 7288 22578 7340 22584
rect 7300 22234 7328 22578
rect 7288 22228 7340 22234
rect 7288 22170 7340 22176
rect 7392 22094 7420 32166
rect 10180 32124 10556 32133
rect 10236 32122 10260 32124
rect 10316 32122 10340 32124
rect 10396 32122 10420 32124
rect 10476 32122 10500 32124
rect 10236 32070 10246 32122
rect 10490 32070 10500 32122
rect 10236 32068 10260 32070
rect 10316 32068 10340 32070
rect 10396 32068 10420 32070
rect 10476 32068 10500 32070
rect 10180 32059 10556 32068
rect 10920 31580 11296 31589
rect 10976 31578 11000 31580
rect 11056 31578 11080 31580
rect 11136 31578 11160 31580
rect 11216 31578 11240 31580
rect 10976 31526 10986 31578
rect 11230 31526 11240 31578
rect 10976 31524 11000 31526
rect 11056 31524 11080 31526
rect 11136 31524 11160 31526
rect 11216 31524 11240 31526
rect 10920 31515 11296 31524
rect 10784 31272 10836 31278
rect 10784 31214 10836 31220
rect 10180 31036 10556 31045
rect 10236 31034 10260 31036
rect 10316 31034 10340 31036
rect 10396 31034 10420 31036
rect 10476 31034 10500 31036
rect 10236 30982 10246 31034
rect 10490 30982 10500 31034
rect 10236 30980 10260 30982
rect 10316 30980 10340 30982
rect 10396 30980 10420 30982
rect 10476 30980 10500 30982
rect 10180 30971 10556 30980
rect 10796 30734 10824 31214
rect 11612 31136 11664 31142
rect 11612 31078 11664 31084
rect 11624 30802 11652 31078
rect 11612 30796 11664 30802
rect 11612 30738 11664 30744
rect 12452 30734 12480 32234
rect 13176 32224 13228 32230
rect 13176 32166 13228 32172
rect 13188 31754 13216 32166
rect 16180 32124 16556 32133
rect 16236 32122 16260 32124
rect 16316 32122 16340 32124
rect 16396 32122 16420 32124
rect 16476 32122 16500 32124
rect 16236 32070 16246 32122
rect 16490 32070 16500 32122
rect 16236 32068 16260 32070
rect 16316 32068 16340 32070
rect 16396 32068 16420 32070
rect 16476 32068 16500 32070
rect 16180 32059 16556 32068
rect 13096 31726 13216 31754
rect 13544 31748 13596 31754
rect 12808 31272 12860 31278
rect 12808 31214 12860 31220
rect 12900 31272 12952 31278
rect 12900 31214 12952 31220
rect 10784 30728 10836 30734
rect 10784 30670 10836 30676
rect 12440 30728 12492 30734
rect 12440 30670 12492 30676
rect 10180 29948 10556 29957
rect 10236 29946 10260 29948
rect 10316 29946 10340 29948
rect 10396 29946 10420 29948
rect 10476 29946 10500 29948
rect 10236 29894 10246 29946
rect 10490 29894 10500 29946
rect 10236 29892 10260 29894
rect 10316 29892 10340 29894
rect 10396 29892 10420 29894
rect 10476 29892 10500 29894
rect 10180 29883 10556 29892
rect 10180 28860 10556 28869
rect 10236 28858 10260 28860
rect 10316 28858 10340 28860
rect 10396 28858 10420 28860
rect 10476 28858 10500 28860
rect 10236 28806 10246 28858
rect 10490 28806 10500 28858
rect 10236 28804 10260 28806
rect 10316 28804 10340 28806
rect 10396 28804 10420 28806
rect 10476 28804 10500 28806
rect 10180 28795 10556 28804
rect 8484 28552 8536 28558
rect 8484 28494 8536 28500
rect 8668 28552 8720 28558
rect 8668 28494 8720 28500
rect 8496 28218 8524 28494
rect 8484 28212 8536 28218
rect 8484 28154 8536 28160
rect 7840 27872 7892 27878
rect 7840 27814 7892 27820
rect 7564 26240 7616 26246
rect 7564 26182 7616 26188
rect 7576 26042 7604 26182
rect 7564 26036 7616 26042
rect 7564 25978 7616 25984
rect 7748 25220 7800 25226
rect 7748 25162 7800 25168
rect 7760 24954 7788 25162
rect 7748 24948 7800 24954
rect 7748 24890 7800 24896
rect 7748 22976 7800 22982
rect 7748 22918 7800 22924
rect 7392 22066 7604 22094
rect 6092 21888 6144 21894
rect 6092 21830 6144 21836
rect 6276 21888 6328 21894
rect 6276 21830 6328 21836
rect 6552 21888 6604 21894
rect 6552 21830 6604 21836
rect 7196 21888 7248 21894
rect 7196 21830 7248 21836
rect 6104 21622 6132 21830
rect 6092 21616 6144 21622
rect 6092 21558 6144 21564
rect 6184 21548 6236 21554
rect 6184 21490 6236 21496
rect 6196 21146 6224 21490
rect 6184 21140 6236 21146
rect 6184 21082 6236 21088
rect 6288 21010 6316 21830
rect 6564 21690 6592 21830
rect 6552 21684 6604 21690
rect 6552 21626 6604 21632
rect 7104 21684 7156 21690
rect 7104 21626 7156 21632
rect 6368 21344 6420 21350
rect 6368 21286 6420 21292
rect 6380 21146 6408 21286
rect 6368 21140 6420 21146
rect 6368 21082 6420 21088
rect 6276 21004 6328 21010
rect 6276 20946 6328 20952
rect 6920 20392 6972 20398
rect 6920 20334 6972 20340
rect 6932 19854 6960 20334
rect 6920 19848 6972 19854
rect 6920 19790 6972 19796
rect 6932 19378 6960 19790
rect 6000 19372 6052 19378
rect 6000 19314 6052 19320
rect 6920 19372 6972 19378
rect 6920 19314 6972 19320
rect 5828 19230 5948 19258
rect 5828 18766 5856 19230
rect 5908 19168 5960 19174
rect 5908 19110 5960 19116
rect 5920 18970 5948 19110
rect 6012 18970 6040 19314
rect 5908 18964 5960 18970
rect 5908 18906 5960 18912
rect 6000 18964 6052 18970
rect 6000 18906 6052 18912
rect 5552 18698 5764 18714
rect 5816 18760 5868 18766
rect 5816 18702 5868 18708
rect 5540 18692 5764 18698
rect 5592 18686 5764 18692
rect 5540 18634 5592 18640
rect 4804 18624 4856 18630
rect 4804 18566 4856 18572
rect 4920 18524 5296 18533
rect 4976 18522 5000 18524
rect 5056 18522 5080 18524
rect 5136 18522 5160 18524
rect 5216 18522 5240 18524
rect 4976 18470 4986 18522
rect 5230 18470 5240 18522
rect 4976 18468 5000 18470
rect 5056 18468 5080 18470
rect 5136 18468 5160 18470
rect 5216 18468 5240 18470
rect 4920 18459 5296 18468
rect 5736 17610 5764 18686
rect 5828 17814 5856 18702
rect 5816 17808 5868 17814
rect 5816 17750 5868 17756
rect 5724 17604 5776 17610
rect 5724 17546 5776 17552
rect 4804 17536 4856 17542
rect 4804 17478 4856 17484
rect 5356 17536 5408 17542
rect 5356 17478 5408 17484
rect 4816 17338 4844 17478
rect 4920 17436 5296 17445
rect 4976 17434 5000 17436
rect 5056 17434 5080 17436
rect 5136 17434 5160 17436
rect 5216 17434 5240 17436
rect 4976 17382 4986 17434
rect 5230 17382 5240 17434
rect 4976 17380 5000 17382
rect 5056 17380 5080 17382
rect 5136 17380 5160 17382
rect 5216 17380 5240 17382
rect 4920 17371 5296 17380
rect 5368 17338 5396 17478
rect 4804 17332 4856 17338
rect 4804 17274 4856 17280
rect 5356 17332 5408 17338
rect 5356 17274 5408 17280
rect 5356 17128 5408 17134
rect 5356 17070 5408 17076
rect 4896 16992 4948 16998
rect 4896 16934 4948 16940
rect 4724 16748 4844 16776
rect 4632 16646 4752 16674
rect 4620 16516 4672 16522
rect 4620 16458 4672 16464
rect 4632 16250 4660 16458
rect 4620 16244 4672 16250
rect 4620 16186 4672 16192
rect 4180 15804 4556 15813
rect 4236 15802 4260 15804
rect 4316 15802 4340 15804
rect 4396 15802 4420 15804
rect 4476 15802 4500 15804
rect 4236 15750 4246 15802
rect 4490 15750 4500 15802
rect 4236 15748 4260 15750
rect 4316 15748 4340 15750
rect 4396 15748 4420 15750
rect 4476 15748 4500 15750
rect 4180 15739 4556 15748
rect 4068 14952 4120 14958
rect 4068 14894 4120 14900
rect 3792 14272 3844 14278
rect 3792 14214 3844 14220
rect 3804 13326 3832 14214
rect 3792 13320 3844 13326
rect 3792 13262 3844 13268
rect 3976 12096 4028 12102
rect 3976 12038 4028 12044
rect 3988 11898 4016 12038
rect 3976 11892 4028 11898
rect 3976 11834 4028 11840
rect 3700 11688 3752 11694
rect 3700 11630 3752 11636
rect 3712 11354 3740 11630
rect 2596 11348 2648 11354
rect 2596 11290 2648 11296
rect 3700 11348 3752 11354
rect 3700 11290 3752 11296
rect 4080 11218 4108 14894
rect 4620 14816 4672 14822
rect 4620 14758 4672 14764
rect 4180 14716 4556 14725
rect 4236 14714 4260 14716
rect 4316 14714 4340 14716
rect 4396 14714 4420 14716
rect 4476 14714 4500 14716
rect 4236 14662 4246 14714
rect 4490 14662 4500 14714
rect 4236 14660 4260 14662
rect 4316 14660 4340 14662
rect 4396 14660 4420 14662
rect 4476 14660 4500 14662
rect 4180 14651 4556 14660
rect 4160 14272 4212 14278
rect 4160 14214 4212 14220
rect 4172 14074 4200 14214
rect 4160 14068 4212 14074
rect 4160 14010 4212 14016
rect 4632 14006 4660 14758
rect 4724 14482 4752 16646
rect 4816 16046 4844 16748
rect 4908 16590 4936 16934
rect 5368 16726 5396 17070
rect 5356 16720 5408 16726
rect 5356 16662 5408 16668
rect 4896 16584 4948 16590
rect 4896 16526 4948 16532
rect 4920 16348 5296 16357
rect 4976 16346 5000 16348
rect 5056 16346 5080 16348
rect 5136 16346 5160 16348
rect 5216 16346 5240 16348
rect 4976 16294 4986 16346
rect 5230 16294 5240 16346
rect 4976 16292 5000 16294
rect 5056 16292 5080 16294
rect 5136 16292 5160 16294
rect 5216 16292 5240 16294
rect 4920 16283 5296 16292
rect 5368 16250 5396 16662
rect 5356 16244 5408 16250
rect 5356 16186 5408 16192
rect 4804 16040 4856 16046
rect 4804 15982 4856 15988
rect 4816 14958 4844 15982
rect 4920 15260 5296 15269
rect 4976 15258 5000 15260
rect 5056 15258 5080 15260
rect 5136 15258 5160 15260
rect 5216 15258 5240 15260
rect 4976 15206 4986 15258
rect 5230 15206 5240 15258
rect 4976 15204 5000 15206
rect 5056 15204 5080 15206
rect 5136 15204 5160 15206
rect 5216 15204 5240 15206
rect 4920 15195 5296 15204
rect 4804 14952 4856 14958
rect 4804 14894 4856 14900
rect 4712 14476 4764 14482
rect 4712 14418 4764 14424
rect 4620 14000 4672 14006
rect 4620 13942 4672 13948
rect 4180 13628 4556 13637
rect 4236 13626 4260 13628
rect 4316 13626 4340 13628
rect 4396 13626 4420 13628
rect 4476 13626 4500 13628
rect 4236 13574 4246 13626
rect 4490 13574 4500 13626
rect 4236 13572 4260 13574
rect 4316 13572 4340 13574
rect 4396 13572 4420 13574
rect 4476 13572 4500 13574
rect 4180 13563 4556 13572
rect 4180 12540 4556 12549
rect 4236 12538 4260 12540
rect 4316 12538 4340 12540
rect 4396 12538 4420 12540
rect 4476 12538 4500 12540
rect 4236 12486 4246 12538
rect 4490 12486 4500 12538
rect 4236 12484 4260 12486
rect 4316 12484 4340 12486
rect 4396 12484 4420 12486
rect 4476 12484 4500 12486
rect 4180 12475 4556 12484
rect 4724 12322 4752 14418
rect 4920 14172 5296 14181
rect 4976 14170 5000 14172
rect 5056 14170 5080 14172
rect 5136 14170 5160 14172
rect 5216 14170 5240 14172
rect 4976 14118 4986 14170
rect 5230 14118 5240 14170
rect 4976 14116 5000 14118
rect 5056 14116 5080 14118
rect 5136 14116 5160 14118
rect 5216 14116 5240 14118
rect 4920 14107 5296 14116
rect 5356 14068 5408 14074
rect 5356 14010 5408 14016
rect 4920 13084 5296 13093
rect 4976 13082 5000 13084
rect 5056 13082 5080 13084
rect 5136 13082 5160 13084
rect 5216 13082 5240 13084
rect 4976 13030 4986 13082
rect 5230 13030 5240 13082
rect 4976 13028 5000 13030
rect 5056 13028 5080 13030
rect 5136 13028 5160 13030
rect 5216 13028 5240 13030
rect 4920 13019 5296 13028
rect 4632 12306 4752 12322
rect 4160 12300 4212 12306
rect 4160 12242 4212 12248
rect 4632 12300 4764 12306
rect 4632 12294 4712 12300
rect 4172 11694 4200 12242
rect 4252 12096 4304 12102
rect 4252 12038 4304 12044
rect 4436 12096 4488 12102
rect 4436 12038 4488 12044
rect 4264 11898 4292 12038
rect 4252 11892 4304 11898
rect 4252 11834 4304 11840
rect 4448 11762 4476 12038
rect 4436 11756 4488 11762
rect 4436 11698 4488 11704
rect 4160 11688 4212 11694
rect 4160 11630 4212 11636
rect 4180 11452 4556 11461
rect 4236 11450 4260 11452
rect 4316 11450 4340 11452
rect 4396 11450 4420 11452
rect 4476 11450 4500 11452
rect 4236 11398 4246 11450
rect 4490 11398 4500 11450
rect 4236 11396 4260 11398
rect 4316 11396 4340 11398
rect 4396 11396 4420 11398
rect 4476 11396 4500 11398
rect 4180 11387 4556 11396
rect 4068 11212 4120 11218
rect 4068 11154 4120 11160
rect 2596 10668 2648 10674
rect 2596 10610 2648 10616
rect 2504 10600 2556 10606
rect 2504 10542 2556 10548
rect 2516 9586 2544 10542
rect 2608 10266 2636 10610
rect 4080 10470 4108 11154
rect 4632 10606 4660 12294
rect 4712 12242 4764 12248
rect 4804 12232 4856 12238
rect 4804 12174 4856 12180
rect 4712 12164 4764 12170
rect 4712 12106 4764 12112
rect 4724 11898 4752 12106
rect 4712 11892 4764 11898
rect 4712 11834 4764 11840
rect 4816 11762 4844 12174
rect 4920 11996 5296 12005
rect 4976 11994 5000 11996
rect 5056 11994 5080 11996
rect 5136 11994 5160 11996
rect 5216 11994 5240 11996
rect 4976 11942 4986 11994
rect 5230 11942 5240 11994
rect 4976 11940 5000 11942
rect 5056 11940 5080 11942
rect 5136 11940 5160 11942
rect 5216 11940 5240 11942
rect 4920 11931 5296 11940
rect 5080 11892 5132 11898
rect 5080 11834 5132 11840
rect 5092 11762 5120 11834
rect 5368 11762 5396 14010
rect 5736 14006 5764 17546
rect 5828 14074 5856 17750
rect 6932 17678 6960 19314
rect 7116 18834 7144 21626
rect 7208 21486 7236 21830
rect 7380 21548 7432 21554
rect 7380 21490 7432 21496
rect 7196 21480 7248 21486
rect 7196 21422 7248 21428
rect 7288 20256 7340 20262
rect 7288 20198 7340 20204
rect 7300 19854 7328 20198
rect 7288 19848 7340 19854
rect 7288 19790 7340 19796
rect 7104 18828 7156 18834
rect 7104 18770 7156 18776
rect 7196 18828 7248 18834
rect 7196 18770 7248 18776
rect 6920 17672 6972 17678
rect 6920 17614 6972 17620
rect 6092 17604 6144 17610
rect 6092 17546 6144 17552
rect 6104 16658 6132 17546
rect 6368 17536 6420 17542
rect 6368 17478 6420 17484
rect 6380 17338 6408 17478
rect 6368 17332 6420 17338
rect 6368 17274 6420 17280
rect 6932 16998 6960 17614
rect 7012 17264 7064 17270
rect 7012 17206 7064 17212
rect 6920 16992 6972 16998
rect 6920 16934 6972 16940
rect 7024 16794 7052 17206
rect 7012 16788 7064 16794
rect 7012 16730 7064 16736
rect 6092 16652 6144 16658
rect 6092 16594 6144 16600
rect 6828 16584 6880 16590
rect 6828 16526 6880 16532
rect 6644 15360 6696 15366
rect 6644 15302 6696 15308
rect 6656 15162 6684 15302
rect 6840 15162 6868 16526
rect 7208 15586 7236 18770
rect 7288 18080 7340 18086
rect 7288 18022 7340 18028
rect 7300 17678 7328 18022
rect 7288 17672 7340 17678
rect 7288 17614 7340 17620
rect 7392 16658 7420 21490
rect 7472 20460 7524 20466
rect 7472 20402 7524 20408
rect 7484 19514 7512 20402
rect 7472 19508 7524 19514
rect 7472 19450 7524 19456
rect 7576 18630 7604 22066
rect 7760 22030 7788 22918
rect 7748 22024 7800 22030
rect 7748 21966 7800 21972
rect 7852 21554 7880 27814
rect 8680 27470 8708 28494
rect 10796 28490 10824 30670
rect 10920 30492 11296 30501
rect 10976 30490 11000 30492
rect 11056 30490 11080 30492
rect 11136 30490 11160 30492
rect 11216 30490 11240 30492
rect 10976 30438 10986 30490
rect 11230 30438 11240 30490
rect 10976 30436 11000 30438
rect 11056 30436 11080 30438
rect 11136 30436 11160 30438
rect 11216 30436 11240 30438
rect 10920 30427 11296 30436
rect 12820 30394 12848 31214
rect 12912 30870 12940 31214
rect 12900 30864 12952 30870
rect 12900 30806 12952 30812
rect 12808 30388 12860 30394
rect 12808 30330 12860 30336
rect 12912 30258 12940 30806
rect 12992 30728 13044 30734
rect 12992 30670 13044 30676
rect 11888 30252 11940 30258
rect 11888 30194 11940 30200
rect 12900 30252 12952 30258
rect 12900 30194 12952 30200
rect 10920 29404 11296 29413
rect 10976 29402 11000 29404
rect 11056 29402 11080 29404
rect 11136 29402 11160 29404
rect 11216 29402 11240 29404
rect 10976 29350 10986 29402
rect 11230 29350 11240 29402
rect 10976 29348 11000 29350
rect 11056 29348 11080 29350
rect 11136 29348 11160 29350
rect 11216 29348 11240 29350
rect 10920 29339 11296 29348
rect 11900 28762 11928 30194
rect 13004 29714 13032 30670
rect 12992 29708 13044 29714
rect 12992 29650 13044 29656
rect 11888 28756 11940 28762
rect 11888 28698 11940 28704
rect 10784 28484 10836 28490
rect 10784 28426 10836 28432
rect 10324 28416 10376 28422
rect 10324 28358 10376 28364
rect 10508 28416 10560 28422
rect 10508 28358 10560 28364
rect 10336 28014 10364 28358
rect 10520 28218 10548 28358
rect 10508 28212 10560 28218
rect 10508 28154 10560 28160
rect 9220 28008 9272 28014
rect 9220 27950 9272 27956
rect 9864 28008 9916 28014
rect 9864 27950 9916 27956
rect 10324 28008 10376 28014
rect 10324 27950 10376 27956
rect 10692 28008 10744 28014
rect 10692 27950 10744 27956
rect 8668 27464 8720 27470
rect 8668 27406 8720 27412
rect 8392 26920 8444 26926
rect 8392 26862 8444 26868
rect 8404 26586 8432 26862
rect 8392 26580 8444 26586
rect 8392 26522 8444 26528
rect 8300 25832 8352 25838
rect 8300 25774 8352 25780
rect 8312 24750 8340 25774
rect 8404 25430 8432 26522
rect 8576 26240 8628 26246
rect 8576 26182 8628 26188
rect 8588 26042 8616 26182
rect 8576 26036 8628 26042
rect 8576 25978 8628 25984
rect 8392 25424 8444 25430
rect 8392 25366 8444 25372
rect 8680 25294 8708 27406
rect 9128 27396 9180 27402
rect 9128 27338 9180 27344
rect 9140 26586 9168 27338
rect 9232 27033 9260 27950
rect 9312 27396 9364 27402
rect 9312 27338 9364 27344
rect 9324 27130 9352 27338
rect 9312 27124 9364 27130
rect 9312 27066 9364 27072
rect 9218 27024 9274 27033
rect 9218 26959 9274 26968
rect 9128 26580 9180 26586
rect 9128 26522 9180 26528
rect 9232 25498 9260 26959
rect 9680 26920 9732 26926
rect 9680 26862 9732 26868
rect 9692 26234 9720 26862
rect 9600 26206 9720 26234
rect 9496 25696 9548 25702
rect 9496 25638 9548 25644
rect 9220 25492 9272 25498
rect 9220 25434 9272 25440
rect 8668 25288 8720 25294
rect 8668 25230 8720 25236
rect 8576 25152 8628 25158
rect 8576 25094 8628 25100
rect 8300 24744 8352 24750
rect 8300 24686 8352 24692
rect 8588 24138 8616 25094
rect 8680 24750 8708 25230
rect 8944 25152 8996 25158
rect 8944 25094 8996 25100
rect 9312 25152 9364 25158
rect 9312 25094 9364 25100
rect 8956 24954 8984 25094
rect 8944 24948 8996 24954
rect 8944 24890 8996 24896
rect 8852 24812 8904 24818
rect 8852 24754 8904 24760
rect 8668 24744 8720 24750
rect 8668 24686 8720 24692
rect 8576 24132 8628 24138
rect 8576 24074 8628 24080
rect 8024 24064 8076 24070
rect 8024 24006 8076 24012
rect 8036 23746 8064 24006
rect 8036 23730 8156 23746
rect 8036 23724 8168 23730
rect 8036 23718 8116 23724
rect 8116 23666 8168 23672
rect 7932 23112 7984 23118
rect 7932 23054 7984 23060
rect 7944 22778 7972 23054
rect 7932 22772 7984 22778
rect 7932 22714 7984 22720
rect 7944 22030 7972 22714
rect 8024 22432 8076 22438
rect 8024 22374 8076 22380
rect 8036 22234 8064 22374
rect 8024 22228 8076 22234
rect 8024 22170 8076 22176
rect 8128 22094 8156 23666
rect 8680 22710 8708 24686
rect 8864 23662 8892 24754
rect 9220 24744 9272 24750
rect 9220 24686 9272 24692
rect 9232 24410 9260 24686
rect 9220 24404 9272 24410
rect 9220 24346 9272 24352
rect 8852 23656 8904 23662
rect 8852 23598 8904 23604
rect 8944 22976 8996 22982
rect 8944 22918 8996 22924
rect 8956 22778 8984 22918
rect 8944 22772 8996 22778
rect 8944 22714 8996 22720
rect 8668 22704 8720 22710
rect 8668 22646 8720 22652
rect 8576 22568 8628 22574
rect 8576 22510 8628 22516
rect 8036 22066 8156 22094
rect 8036 22030 8064 22066
rect 7932 22024 7984 22030
rect 7932 21966 7984 21972
rect 8024 22024 8076 22030
rect 8024 21966 8076 21972
rect 8484 21888 8536 21894
rect 8484 21830 8536 21836
rect 8206 21584 8262 21593
rect 7840 21548 7892 21554
rect 8206 21519 8208 21528
rect 7840 21490 7892 21496
rect 8260 21519 8262 21528
rect 8208 21490 8260 21496
rect 8220 20754 8248 21490
rect 8496 20942 8524 21830
rect 8484 20936 8536 20942
rect 8484 20878 8536 20884
rect 8392 20868 8444 20874
rect 8392 20810 8444 20816
rect 8220 20726 8340 20754
rect 8312 20534 8340 20726
rect 8300 20528 8352 20534
rect 8300 20470 8352 20476
rect 7748 20460 7800 20466
rect 7748 20402 7800 20408
rect 7760 19242 7788 20402
rect 8404 20346 8432 20810
rect 8312 20318 8432 20346
rect 8312 19310 8340 20318
rect 8208 19304 8260 19310
rect 8208 19246 8260 19252
rect 8300 19304 8352 19310
rect 8300 19246 8352 19252
rect 7748 19236 7800 19242
rect 7748 19178 7800 19184
rect 7760 18834 7788 19178
rect 7748 18828 7800 18834
rect 7748 18770 7800 18776
rect 7564 18624 7616 18630
rect 7564 18566 7616 18572
rect 8116 18216 8168 18222
rect 8116 18158 8168 18164
rect 7840 16992 7892 16998
rect 7840 16934 7892 16940
rect 8024 16992 8076 16998
rect 8024 16934 8076 16940
rect 7852 16658 7880 16934
rect 7380 16652 7432 16658
rect 7380 16594 7432 16600
rect 7840 16652 7892 16658
rect 7840 16594 7892 16600
rect 8036 16590 8064 16934
rect 8024 16584 8076 16590
rect 8024 16526 8076 16532
rect 7116 15558 7236 15586
rect 6644 15156 6696 15162
rect 6644 15098 6696 15104
rect 6828 15156 6880 15162
rect 6828 15098 6880 15104
rect 7116 14958 7144 15558
rect 7196 15496 7248 15502
rect 7196 15438 7248 15444
rect 7840 15496 7892 15502
rect 7840 15438 7892 15444
rect 7104 14952 7156 14958
rect 7104 14894 7156 14900
rect 6368 14816 6420 14822
rect 6368 14758 6420 14764
rect 6000 14340 6052 14346
rect 6000 14282 6052 14288
rect 6012 14074 6040 14282
rect 6380 14074 6408 14758
rect 7208 14618 7236 15438
rect 7564 14816 7616 14822
rect 7564 14758 7616 14764
rect 7196 14612 7248 14618
rect 7196 14554 7248 14560
rect 7012 14340 7064 14346
rect 7012 14282 7064 14288
rect 7024 14074 7052 14282
rect 7576 14074 7604 14758
rect 7852 14618 7880 15438
rect 8128 15162 8156 18158
rect 8220 18154 8248 19246
rect 8588 18306 8616 22510
rect 8680 21622 8708 22646
rect 8944 22024 8996 22030
rect 8944 21966 8996 21972
rect 8668 21616 8720 21622
rect 8668 21558 8720 21564
rect 8760 21616 8812 21622
rect 8760 21558 8812 21564
rect 8772 20806 8800 21558
rect 8852 21548 8904 21554
rect 8852 21490 8904 21496
rect 8760 20800 8812 20806
rect 8760 20742 8812 20748
rect 8772 20466 8800 20742
rect 8760 20460 8812 20466
rect 8760 20402 8812 20408
rect 8864 20398 8892 21490
rect 8956 21146 8984 21966
rect 9220 21956 9272 21962
rect 9220 21898 9272 21904
rect 8944 21140 8996 21146
rect 8944 21082 8996 21088
rect 9232 20874 9260 21898
rect 9324 21842 9352 25094
rect 9508 24410 9536 25638
rect 9600 25378 9628 26206
rect 9876 25906 9904 27950
rect 10180 27772 10556 27781
rect 10236 27770 10260 27772
rect 10316 27770 10340 27772
rect 10396 27770 10420 27772
rect 10476 27770 10500 27772
rect 10236 27718 10246 27770
rect 10490 27718 10500 27770
rect 10236 27716 10260 27718
rect 10316 27716 10340 27718
rect 10396 27716 10420 27718
rect 10476 27716 10500 27718
rect 10180 27707 10556 27716
rect 10600 27396 10652 27402
rect 10600 27338 10652 27344
rect 10048 27328 10100 27334
rect 10048 27270 10100 27276
rect 10508 27328 10560 27334
rect 10508 27270 10560 27276
rect 9956 26444 10008 26450
rect 9956 26386 10008 26392
rect 9680 25900 9732 25906
rect 9680 25842 9732 25848
rect 9864 25900 9916 25906
rect 9864 25842 9916 25848
rect 9692 25498 9720 25842
rect 9680 25492 9732 25498
rect 9680 25434 9732 25440
rect 9864 25424 9916 25430
rect 9600 25350 9720 25378
rect 9864 25366 9916 25372
rect 9692 24614 9720 25350
rect 9772 25152 9824 25158
rect 9772 25094 9824 25100
rect 9680 24608 9732 24614
rect 9680 24550 9732 24556
rect 9496 24404 9548 24410
rect 9496 24346 9548 24352
rect 9404 23316 9456 23322
rect 9404 23258 9456 23264
rect 9416 22642 9444 23258
rect 9404 22636 9456 22642
rect 9404 22578 9456 22584
rect 9416 21962 9444 22578
rect 9404 21956 9456 21962
rect 9404 21898 9456 21904
rect 9324 21814 9444 21842
rect 9416 21400 9444 21814
rect 9508 21554 9536 24346
rect 9784 23882 9812 25094
rect 9692 23854 9812 23882
rect 9588 23656 9640 23662
rect 9588 23598 9640 23604
rect 9600 22574 9628 23598
rect 9588 22568 9640 22574
rect 9588 22510 9640 22516
rect 9588 22092 9640 22098
rect 9588 22034 9640 22040
rect 9600 21690 9628 22034
rect 9588 21684 9640 21690
rect 9588 21626 9640 21632
rect 9496 21548 9548 21554
rect 9496 21490 9548 21496
rect 9416 21372 9536 21400
rect 9312 21344 9364 21350
rect 9364 21292 9444 21298
rect 9312 21286 9444 21292
rect 9324 21270 9444 21286
rect 9220 20868 9272 20874
rect 9220 20810 9272 20816
rect 9312 20800 9364 20806
rect 9312 20742 9364 20748
rect 9324 20602 9352 20742
rect 9312 20596 9364 20602
rect 9312 20538 9364 20544
rect 8852 20392 8904 20398
rect 8852 20334 8904 20340
rect 9416 19802 9444 21270
rect 9508 20466 9536 21372
rect 9692 21010 9720 23854
rect 9772 23792 9824 23798
rect 9772 23734 9824 23740
rect 9680 21004 9732 21010
rect 9680 20946 9732 20952
rect 9784 20466 9812 23734
rect 9876 23526 9904 25366
rect 9968 25294 9996 26386
rect 10060 25906 10088 27270
rect 10520 27130 10548 27270
rect 10508 27124 10560 27130
rect 10508 27066 10560 27072
rect 10612 26926 10640 27338
rect 10600 26920 10652 26926
rect 10600 26862 10652 26868
rect 10180 26684 10556 26693
rect 10236 26682 10260 26684
rect 10316 26682 10340 26684
rect 10396 26682 10420 26684
rect 10476 26682 10500 26684
rect 10236 26630 10246 26682
rect 10490 26630 10500 26682
rect 10236 26628 10260 26630
rect 10316 26628 10340 26630
rect 10396 26628 10420 26630
rect 10476 26628 10500 26630
rect 10180 26619 10556 26628
rect 10048 25900 10100 25906
rect 10048 25842 10100 25848
rect 10140 25900 10192 25906
rect 10140 25842 10192 25848
rect 10152 25702 10180 25842
rect 10140 25696 10192 25702
rect 10140 25638 10192 25644
rect 10180 25596 10556 25605
rect 10236 25594 10260 25596
rect 10316 25594 10340 25596
rect 10396 25594 10420 25596
rect 10476 25594 10500 25596
rect 10236 25542 10246 25594
rect 10490 25542 10500 25594
rect 10236 25540 10260 25542
rect 10316 25540 10340 25542
rect 10396 25540 10420 25542
rect 10476 25540 10500 25542
rect 10180 25531 10556 25540
rect 9956 25288 10008 25294
rect 9956 25230 10008 25236
rect 10048 25220 10100 25226
rect 10048 25162 10100 25168
rect 9956 24064 10008 24070
rect 9956 24006 10008 24012
rect 9864 23520 9916 23526
rect 9864 23462 9916 23468
rect 9864 23044 9916 23050
rect 9864 22986 9916 22992
rect 9876 22778 9904 22986
rect 9864 22772 9916 22778
rect 9864 22714 9916 22720
rect 9864 22568 9916 22574
rect 9864 22510 9916 22516
rect 9876 21486 9904 22510
rect 9968 22250 9996 24006
rect 10060 23798 10088 25162
rect 10612 25158 10640 26862
rect 10704 25906 10732 27950
rect 10692 25900 10744 25906
rect 10692 25842 10744 25848
rect 10704 25430 10732 25842
rect 10692 25424 10744 25430
rect 10692 25366 10744 25372
rect 10796 25294 10824 28426
rect 10920 28316 11296 28325
rect 10976 28314 11000 28316
rect 11056 28314 11080 28316
rect 11136 28314 11160 28316
rect 11216 28314 11240 28316
rect 10976 28262 10986 28314
rect 11230 28262 11240 28314
rect 10976 28260 11000 28262
rect 11056 28260 11080 28262
rect 11136 28260 11160 28262
rect 11216 28260 11240 28262
rect 10920 28251 11296 28260
rect 11900 28082 11928 28698
rect 11888 28076 11940 28082
rect 11888 28018 11940 28024
rect 11336 27872 11388 27878
rect 11336 27814 11388 27820
rect 10920 27228 11296 27237
rect 10976 27226 11000 27228
rect 11056 27226 11080 27228
rect 11136 27226 11160 27228
rect 11216 27226 11240 27228
rect 10976 27174 10986 27226
rect 11230 27174 11240 27226
rect 10976 27172 11000 27174
rect 11056 27172 11080 27174
rect 11136 27172 11160 27174
rect 11216 27172 11240 27174
rect 10920 27163 11296 27172
rect 11348 27062 11376 27814
rect 11336 27056 11388 27062
rect 11336 26998 11388 27004
rect 12532 26920 12584 26926
rect 12532 26862 12584 26868
rect 11336 26240 11388 26246
rect 11336 26182 11388 26188
rect 10920 26140 11296 26149
rect 10976 26138 11000 26140
rect 11056 26138 11080 26140
rect 11136 26138 11160 26140
rect 11216 26138 11240 26140
rect 10976 26086 10986 26138
rect 11230 26086 11240 26138
rect 10976 26084 11000 26086
rect 11056 26084 11080 26086
rect 11136 26084 11160 26086
rect 11216 26084 11240 26086
rect 10920 26075 11296 26084
rect 11348 25770 11376 26182
rect 11336 25764 11388 25770
rect 11336 25706 11388 25712
rect 11612 25764 11664 25770
rect 11612 25706 11664 25712
rect 11428 25696 11480 25702
rect 11428 25638 11480 25644
rect 10784 25288 10836 25294
rect 10784 25230 10836 25236
rect 10600 25152 10652 25158
rect 10600 25094 10652 25100
rect 10690 24712 10746 24721
rect 10600 24676 10652 24682
rect 10690 24647 10692 24656
rect 10600 24618 10652 24624
rect 10744 24647 10746 24656
rect 10692 24618 10744 24624
rect 10180 24508 10556 24517
rect 10236 24506 10260 24508
rect 10316 24506 10340 24508
rect 10396 24506 10420 24508
rect 10476 24506 10500 24508
rect 10236 24454 10246 24506
rect 10490 24454 10500 24506
rect 10236 24452 10260 24454
rect 10316 24452 10340 24454
rect 10396 24452 10420 24454
rect 10476 24452 10500 24454
rect 10180 24443 10556 24452
rect 10048 23792 10100 23798
rect 10048 23734 10100 23740
rect 10048 23520 10100 23526
rect 10048 23462 10100 23468
rect 10060 22574 10088 23462
rect 10180 23420 10556 23429
rect 10236 23418 10260 23420
rect 10316 23418 10340 23420
rect 10396 23418 10420 23420
rect 10476 23418 10500 23420
rect 10236 23366 10246 23418
rect 10490 23366 10500 23418
rect 10236 23364 10260 23366
rect 10316 23364 10340 23366
rect 10396 23364 10420 23366
rect 10476 23364 10500 23366
rect 10180 23355 10556 23364
rect 10048 22568 10100 22574
rect 10048 22510 10100 22516
rect 10180 22332 10556 22341
rect 10236 22330 10260 22332
rect 10316 22330 10340 22332
rect 10396 22330 10420 22332
rect 10476 22330 10500 22332
rect 10236 22278 10246 22330
rect 10490 22278 10500 22330
rect 10236 22276 10260 22278
rect 10316 22276 10340 22278
rect 10396 22276 10420 22278
rect 10476 22276 10500 22278
rect 10180 22267 10556 22276
rect 9968 22222 10088 22250
rect 10060 22216 10088 22222
rect 10140 22228 10192 22234
rect 10060 22188 10140 22216
rect 10140 22170 10192 22176
rect 10232 22160 10284 22166
rect 10612 22114 10640 24618
rect 10704 24206 10732 24618
rect 10692 24200 10744 24206
rect 10692 24142 10744 24148
rect 10692 24064 10744 24070
rect 10692 24006 10744 24012
rect 10232 22102 10284 22108
rect 10048 21548 10100 21554
rect 10244 21536 10272 22102
rect 10520 22086 10640 22114
rect 10416 21888 10468 21894
rect 10416 21830 10468 21836
rect 10428 21622 10456 21830
rect 10416 21616 10468 21622
rect 10416 21558 10468 21564
rect 10100 21508 10272 21536
rect 10048 21490 10100 21496
rect 9864 21480 9916 21486
rect 9864 21422 9916 21428
rect 10520 21400 10548 22086
rect 10600 22024 10652 22030
rect 10600 21966 10652 21972
rect 10060 21372 10548 21400
rect 10060 21078 10088 21372
rect 10180 21244 10556 21253
rect 10236 21242 10260 21244
rect 10316 21242 10340 21244
rect 10396 21242 10420 21244
rect 10476 21242 10500 21244
rect 10236 21190 10246 21242
rect 10490 21190 10500 21242
rect 10236 21188 10260 21190
rect 10316 21188 10340 21190
rect 10396 21188 10420 21190
rect 10476 21188 10500 21190
rect 10180 21179 10556 21188
rect 10612 21146 10640 21966
rect 10704 21350 10732 24006
rect 10796 22166 10824 25230
rect 11336 25220 11388 25226
rect 11336 25162 11388 25168
rect 10920 25052 11296 25061
rect 10976 25050 11000 25052
rect 11056 25050 11080 25052
rect 11136 25050 11160 25052
rect 11216 25050 11240 25052
rect 10976 24998 10986 25050
rect 11230 24998 11240 25050
rect 10976 24996 11000 24998
rect 11056 24996 11080 24998
rect 11136 24996 11160 24998
rect 11216 24996 11240 24998
rect 10920 24987 11296 24996
rect 11348 24954 11376 25162
rect 11336 24948 11388 24954
rect 11336 24890 11388 24896
rect 11440 24206 11468 25638
rect 11428 24200 11480 24206
rect 11428 24142 11480 24148
rect 10920 23964 11296 23973
rect 10976 23962 11000 23964
rect 11056 23962 11080 23964
rect 11136 23962 11160 23964
rect 11216 23962 11240 23964
rect 10976 23910 10986 23962
rect 11230 23910 11240 23962
rect 10976 23908 11000 23910
rect 11056 23908 11080 23910
rect 11136 23908 11160 23910
rect 11216 23908 11240 23910
rect 10920 23899 11296 23908
rect 10920 22876 11296 22885
rect 10976 22874 11000 22876
rect 11056 22874 11080 22876
rect 11136 22874 11160 22876
rect 11216 22874 11240 22876
rect 10976 22822 10986 22874
rect 11230 22822 11240 22874
rect 10976 22820 11000 22822
rect 11056 22820 11080 22822
rect 11136 22820 11160 22822
rect 11216 22820 11240 22822
rect 10920 22811 11296 22820
rect 11060 22432 11112 22438
rect 11060 22374 11112 22380
rect 10784 22160 10836 22166
rect 10784 22102 10836 22108
rect 11072 22030 11100 22374
rect 11060 22024 11112 22030
rect 11060 21966 11112 21972
rect 10784 21956 10836 21962
rect 10784 21898 10836 21904
rect 11336 21956 11388 21962
rect 11336 21898 11388 21904
rect 10796 21690 10824 21898
rect 10920 21788 11296 21797
rect 10976 21786 11000 21788
rect 11056 21786 11080 21788
rect 11136 21786 11160 21788
rect 11216 21786 11240 21788
rect 10976 21734 10986 21786
rect 11230 21734 11240 21786
rect 10976 21732 11000 21734
rect 11056 21732 11080 21734
rect 11136 21732 11160 21734
rect 11216 21732 11240 21734
rect 10920 21723 11296 21732
rect 10784 21684 10836 21690
rect 10784 21626 10836 21632
rect 11348 21593 11376 21898
rect 11334 21584 11390 21593
rect 11334 21519 11390 21528
rect 10692 21344 10744 21350
rect 10692 21286 10744 21292
rect 10600 21140 10652 21146
rect 10600 21082 10652 21088
rect 10048 21072 10100 21078
rect 10048 21014 10100 21020
rect 9864 20936 9916 20942
rect 9864 20878 9916 20884
rect 9496 20460 9548 20466
rect 9496 20402 9548 20408
rect 9772 20460 9824 20466
rect 9772 20402 9824 20408
rect 9508 20346 9536 20402
rect 9508 20330 9812 20346
rect 9508 20324 9824 20330
rect 9508 20318 9772 20324
rect 9772 20266 9824 20272
rect 9496 20256 9548 20262
rect 9496 20198 9548 20204
rect 9508 19922 9536 20198
rect 9496 19916 9548 19922
rect 9496 19858 9548 19864
rect 9416 19774 9536 19802
rect 8944 19712 8996 19718
rect 8944 19654 8996 19660
rect 8956 19514 8984 19654
rect 8944 19508 8996 19514
rect 8944 19450 8996 19456
rect 8496 18278 8616 18306
rect 8496 18222 8524 18278
rect 8484 18216 8536 18222
rect 8484 18158 8536 18164
rect 9220 18216 9272 18222
rect 9220 18158 9272 18164
rect 8208 18148 8260 18154
rect 8208 18090 8260 18096
rect 8116 15156 8168 15162
rect 8116 15098 8168 15104
rect 7932 15020 7984 15026
rect 7932 14962 7984 14968
rect 7944 14618 7972 14962
rect 8220 14958 8248 18090
rect 8300 15496 8352 15502
rect 8300 15438 8352 15444
rect 8208 14952 8260 14958
rect 8208 14894 8260 14900
rect 7840 14612 7892 14618
rect 7840 14554 7892 14560
rect 7932 14612 7984 14618
rect 7932 14554 7984 14560
rect 7852 14346 7880 14554
rect 8312 14414 8340 15438
rect 8300 14408 8352 14414
rect 8300 14350 8352 14356
rect 7840 14340 7892 14346
rect 7840 14282 7892 14288
rect 5816 14068 5868 14074
rect 5816 14010 5868 14016
rect 6000 14068 6052 14074
rect 6000 14010 6052 14016
rect 6368 14068 6420 14074
rect 6368 14010 6420 14016
rect 7012 14068 7064 14074
rect 7012 14010 7064 14016
rect 7564 14068 7616 14074
rect 7564 14010 7616 14016
rect 5448 14000 5500 14006
rect 5448 13942 5500 13948
rect 5724 14000 5776 14006
rect 5724 13942 5776 13948
rect 5460 12374 5488 13942
rect 8312 12850 8340 14350
rect 8300 12844 8352 12850
rect 8300 12786 8352 12792
rect 5448 12368 5500 12374
rect 5448 12310 5500 12316
rect 5460 11898 5488 12310
rect 7196 12300 7248 12306
rect 7196 12242 7248 12248
rect 7012 12232 7064 12238
rect 7012 12174 7064 12180
rect 6368 12096 6420 12102
rect 6368 12038 6420 12044
rect 6828 12096 6880 12102
rect 6828 12038 6880 12044
rect 6920 12096 6972 12102
rect 6920 12038 6972 12044
rect 6380 11898 6408 12038
rect 6840 11898 6868 12038
rect 5448 11892 5500 11898
rect 5448 11834 5500 11840
rect 6368 11892 6420 11898
rect 6368 11834 6420 11840
rect 6828 11892 6880 11898
rect 6828 11834 6880 11840
rect 4804 11756 4856 11762
rect 4804 11698 4856 11704
rect 5080 11756 5132 11762
rect 5080 11698 5132 11704
rect 5172 11756 5224 11762
rect 5172 11698 5224 11704
rect 5356 11756 5408 11762
rect 5356 11698 5408 11704
rect 5184 11150 5212 11698
rect 5172 11144 5224 11150
rect 5172 11086 5224 11092
rect 5460 11098 5488 11834
rect 6184 11756 6236 11762
rect 6184 11698 6236 11704
rect 6368 11756 6420 11762
rect 6368 11698 6420 11704
rect 5632 11688 5684 11694
rect 5632 11630 5684 11636
rect 5644 11354 5672 11630
rect 6196 11354 6224 11698
rect 5632 11348 5684 11354
rect 5632 11290 5684 11296
rect 6184 11348 6236 11354
rect 6184 11290 6236 11296
rect 5908 11212 5960 11218
rect 5908 11154 5960 11160
rect 5460 11070 5672 11098
rect 4920 10908 5296 10917
rect 4976 10906 5000 10908
rect 5056 10906 5080 10908
rect 5136 10906 5160 10908
rect 5216 10906 5240 10908
rect 4976 10854 4986 10906
rect 5230 10854 5240 10906
rect 4976 10852 5000 10854
rect 5056 10852 5080 10854
rect 5136 10852 5160 10854
rect 5216 10852 5240 10854
rect 4920 10843 5296 10852
rect 4712 10736 4764 10742
rect 4712 10678 4764 10684
rect 4620 10600 4672 10606
rect 4620 10542 4672 10548
rect 3976 10464 4028 10470
rect 3976 10406 4028 10412
rect 4068 10464 4120 10470
rect 4724 10418 4752 10678
rect 5644 10674 5672 11070
rect 5172 10668 5224 10674
rect 5172 10610 5224 10616
rect 5632 10668 5684 10674
rect 5632 10610 5684 10616
rect 4068 10406 4120 10412
rect 3988 10266 4016 10406
rect 2596 10260 2648 10266
rect 2596 10202 2648 10208
rect 3976 10260 4028 10266
rect 3976 10202 4028 10208
rect 4080 10130 4108 10406
rect 4632 10390 4752 10418
rect 4180 10364 4556 10373
rect 4236 10362 4260 10364
rect 4316 10362 4340 10364
rect 4396 10362 4420 10364
rect 4476 10362 4500 10364
rect 4236 10310 4246 10362
rect 4490 10310 4500 10362
rect 4236 10308 4260 10310
rect 4316 10308 4340 10310
rect 4396 10308 4420 10310
rect 4476 10308 4500 10310
rect 4180 10299 4556 10308
rect 4068 10124 4120 10130
rect 4068 10066 4120 10072
rect 3792 9920 3844 9926
rect 3792 9862 3844 9868
rect 4528 9920 4580 9926
rect 4632 9874 4660 10390
rect 5184 10062 5212 10610
rect 4712 10056 4764 10062
rect 4712 9998 4764 10004
rect 5172 10056 5224 10062
rect 5172 9998 5224 10004
rect 4580 9868 4660 9874
rect 4528 9862 4660 9868
rect 2504 9580 2556 9586
rect 2504 9522 2556 9528
rect 2780 9580 2832 9586
rect 2780 9522 2832 9528
rect 2516 7954 2544 9522
rect 2792 9178 2820 9522
rect 2780 9172 2832 9178
rect 2780 9114 2832 9120
rect 3804 8974 3832 9862
rect 4540 9846 4660 9862
rect 4180 9276 4556 9285
rect 4236 9274 4260 9276
rect 4316 9274 4340 9276
rect 4396 9274 4420 9276
rect 4476 9274 4500 9276
rect 4236 9222 4246 9274
rect 4490 9222 4500 9274
rect 4236 9220 4260 9222
rect 4316 9220 4340 9222
rect 4396 9220 4420 9222
rect 4476 9220 4500 9222
rect 4180 9211 4556 9220
rect 3792 8968 3844 8974
rect 3792 8910 3844 8916
rect 4180 8188 4556 8197
rect 4236 8186 4260 8188
rect 4316 8186 4340 8188
rect 4396 8186 4420 8188
rect 4476 8186 4500 8188
rect 4236 8134 4246 8186
rect 4490 8134 4500 8186
rect 4236 8132 4260 8134
rect 4316 8132 4340 8134
rect 4396 8132 4420 8134
rect 4476 8132 4500 8134
rect 4180 8123 4556 8132
rect 2504 7948 2556 7954
rect 2504 7890 2556 7896
rect 4180 7100 4556 7109
rect 4236 7098 4260 7100
rect 4316 7098 4340 7100
rect 4396 7098 4420 7100
rect 4476 7098 4500 7100
rect 4236 7046 4246 7098
rect 4490 7046 4500 7098
rect 4236 7044 4260 7046
rect 4316 7044 4340 7046
rect 4396 7044 4420 7046
rect 4476 7044 4500 7046
rect 4180 7035 4556 7044
rect 4632 6458 4660 9846
rect 4724 9450 4752 9998
rect 4920 9820 5296 9829
rect 4976 9818 5000 9820
rect 5056 9818 5080 9820
rect 5136 9818 5160 9820
rect 5216 9818 5240 9820
rect 4976 9766 4986 9818
rect 5230 9766 5240 9818
rect 4976 9764 5000 9766
rect 5056 9764 5080 9766
rect 5136 9764 5160 9766
rect 5216 9764 5240 9766
rect 4920 9755 5296 9764
rect 4712 9444 4764 9450
rect 4712 9386 4764 9392
rect 4920 8732 5296 8741
rect 4976 8730 5000 8732
rect 5056 8730 5080 8732
rect 5136 8730 5160 8732
rect 5216 8730 5240 8732
rect 4976 8678 4986 8730
rect 5230 8678 5240 8730
rect 4976 8676 5000 8678
rect 5056 8676 5080 8678
rect 5136 8676 5160 8678
rect 5216 8676 5240 8678
rect 4920 8667 5296 8676
rect 5816 8356 5868 8362
rect 5816 8298 5868 8304
rect 5356 7880 5408 7886
rect 5356 7822 5408 7828
rect 4920 7644 5296 7653
rect 4976 7642 5000 7644
rect 5056 7642 5080 7644
rect 5136 7642 5160 7644
rect 5216 7642 5240 7644
rect 4976 7590 4986 7642
rect 5230 7590 5240 7642
rect 4976 7588 5000 7590
rect 5056 7588 5080 7590
rect 5136 7588 5160 7590
rect 5216 7588 5240 7590
rect 4920 7579 5296 7588
rect 5368 6866 5396 7822
rect 5632 7812 5684 7818
rect 5632 7754 5684 7760
rect 5644 7546 5672 7754
rect 5632 7540 5684 7546
rect 5632 7482 5684 7488
rect 5356 6860 5408 6866
rect 5408 6820 5488 6848
rect 5356 6802 5408 6808
rect 4920 6556 5296 6565
rect 4976 6554 5000 6556
rect 5056 6554 5080 6556
rect 5136 6554 5160 6556
rect 5216 6554 5240 6556
rect 4976 6502 4986 6554
rect 5230 6502 5240 6554
rect 4976 6500 5000 6502
rect 5056 6500 5080 6502
rect 5136 6500 5160 6502
rect 5216 6500 5240 6502
rect 4920 6491 5296 6500
rect 4620 6452 4672 6458
rect 4620 6394 4672 6400
rect 5356 6452 5408 6458
rect 5356 6394 5408 6400
rect 940 6316 992 6322
rect 940 6258 992 6264
rect 952 6225 980 6258
rect 938 6216 994 6225
rect 938 6151 994 6160
rect 4180 6012 4556 6021
rect 4236 6010 4260 6012
rect 4316 6010 4340 6012
rect 4396 6010 4420 6012
rect 4476 6010 4500 6012
rect 4236 5958 4246 6010
rect 4490 5958 4500 6010
rect 4236 5956 4260 5958
rect 4316 5956 4340 5958
rect 4396 5956 4420 5958
rect 4476 5956 4500 5958
rect 4180 5947 4556 5956
rect 5368 5642 5396 6394
rect 5460 6322 5488 6820
rect 5828 6730 5856 8298
rect 5920 7478 5948 11154
rect 6196 10606 6224 11290
rect 6380 11150 6408 11698
rect 6736 11552 6788 11558
rect 6736 11494 6788 11500
rect 6368 11144 6420 11150
rect 6368 11086 6420 11092
rect 6748 10606 6776 11494
rect 6932 10810 6960 12038
rect 7024 10810 7052 12174
rect 7104 12164 7156 12170
rect 7104 12106 7156 12112
rect 7116 11150 7144 12106
rect 7104 11144 7156 11150
rect 7104 11086 7156 11092
rect 6920 10804 6972 10810
rect 6920 10746 6972 10752
rect 7012 10804 7064 10810
rect 7012 10746 7064 10752
rect 7208 10742 7236 12242
rect 8024 12232 8076 12238
rect 8496 12186 8524 18158
rect 9232 17882 9260 18158
rect 9508 18086 9536 19774
rect 9876 19378 9904 20878
rect 9864 19372 9916 19378
rect 9864 19314 9916 19320
rect 10060 19258 10088 21014
rect 10180 20156 10556 20165
rect 10236 20154 10260 20156
rect 10316 20154 10340 20156
rect 10396 20154 10420 20156
rect 10476 20154 10500 20156
rect 10236 20102 10246 20154
rect 10490 20102 10500 20154
rect 10236 20100 10260 20102
rect 10316 20100 10340 20102
rect 10396 20100 10420 20102
rect 10476 20100 10500 20102
rect 10180 20091 10556 20100
rect 10600 19372 10652 19378
rect 10600 19314 10652 19320
rect 9784 19230 10088 19258
rect 9496 18080 9548 18086
rect 9496 18022 9548 18028
rect 8852 17876 8904 17882
rect 8852 17818 8904 17824
rect 9220 17876 9272 17882
rect 9220 17818 9272 17824
rect 8864 17270 8892 17818
rect 8852 17264 8904 17270
rect 8852 17206 8904 17212
rect 8760 17196 8812 17202
rect 8760 17138 8812 17144
rect 8772 16794 8800 17138
rect 9128 17060 9180 17066
rect 9128 17002 9180 17008
rect 9036 16992 9088 16998
rect 9036 16934 9088 16940
rect 8760 16788 8812 16794
rect 8760 16730 8812 16736
rect 9048 16114 9076 16934
rect 9140 16726 9168 17002
rect 9128 16720 9180 16726
rect 9128 16662 9180 16668
rect 9508 16250 9536 18022
rect 9680 16992 9732 16998
rect 9680 16934 9732 16940
rect 9588 16448 9640 16454
rect 9588 16390 9640 16396
rect 9496 16244 9548 16250
rect 9496 16186 9548 16192
rect 9600 16114 9628 16390
rect 9692 16114 9720 16934
rect 8944 16108 8996 16114
rect 8944 16050 8996 16056
rect 9036 16108 9088 16114
rect 9036 16050 9088 16056
rect 9312 16108 9364 16114
rect 9312 16050 9364 16056
rect 9588 16108 9640 16114
rect 9588 16050 9640 16056
rect 9680 16108 9732 16114
rect 9680 16050 9732 16056
rect 8956 15706 8984 16050
rect 9324 15706 9352 16050
rect 9784 15994 9812 19230
rect 10180 19068 10556 19077
rect 10236 19066 10260 19068
rect 10316 19066 10340 19068
rect 10396 19066 10420 19068
rect 10476 19066 10500 19068
rect 10236 19014 10246 19066
rect 10490 19014 10500 19066
rect 10236 19012 10260 19014
rect 10316 19012 10340 19014
rect 10396 19012 10420 19014
rect 10476 19012 10500 19014
rect 10180 19003 10556 19012
rect 10612 18970 10640 19314
rect 10600 18964 10652 18970
rect 10600 18906 10652 18912
rect 10704 18578 10732 21286
rect 10968 21072 11020 21078
rect 11020 21020 11284 21026
rect 10968 21014 11284 21020
rect 10876 21004 10928 21010
rect 10980 20998 11284 21014
rect 10876 20946 10928 20952
rect 10888 20806 10916 20946
rect 11256 20942 11284 20998
rect 11348 20942 11376 21519
rect 11520 21344 11572 21350
rect 11520 21286 11572 21292
rect 11532 21078 11560 21286
rect 11520 21072 11572 21078
rect 11520 21014 11572 21020
rect 11428 21004 11480 21010
rect 11428 20946 11480 20952
rect 11244 20936 11296 20942
rect 11244 20878 11296 20884
rect 11336 20936 11388 20942
rect 11336 20878 11388 20884
rect 10876 20800 10928 20806
rect 10876 20742 10928 20748
rect 10920 20700 11296 20709
rect 10976 20698 11000 20700
rect 11056 20698 11080 20700
rect 11136 20698 11160 20700
rect 11216 20698 11240 20700
rect 10976 20646 10986 20698
rect 11230 20646 11240 20698
rect 10976 20644 11000 20646
rect 11056 20644 11080 20646
rect 11136 20644 11160 20646
rect 11216 20644 11240 20646
rect 10920 20635 11296 20644
rect 11440 20602 11468 20946
rect 10784 20596 10836 20602
rect 10784 20538 10836 20544
rect 11428 20596 11480 20602
rect 11428 20538 11480 20544
rect 9692 15966 9812 15994
rect 9968 18550 10732 18578
rect 8944 15700 8996 15706
rect 8944 15642 8996 15648
rect 9312 15700 9364 15706
rect 9312 15642 9364 15648
rect 8760 15632 8812 15638
rect 8760 15574 8812 15580
rect 8576 15496 8628 15502
rect 8576 15438 8628 15444
rect 8588 15162 8616 15438
rect 8772 15434 8800 15574
rect 8760 15428 8812 15434
rect 8760 15370 8812 15376
rect 8576 15156 8628 15162
rect 8576 15098 8628 15104
rect 9036 12912 9088 12918
rect 9036 12854 9088 12860
rect 8944 12776 8996 12782
rect 8944 12718 8996 12724
rect 8956 12442 8984 12718
rect 8944 12436 8996 12442
rect 8944 12378 8996 12384
rect 8024 12174 8076 12180
rect 7932 12096 7984 12102
rect 7932 12038 7984 12044
rect 7944 11762 7972 12038
rect 8036 11898 8064 12174
rect 8404 12158 8524 12186
rect 8668 12232 8720 12238
rect 8668 12174 8720 12180
rect 8024 11892 8076 11898
rect 8024 11834 8076 11840
rect 7932 11756 7984 11762
rect 7932 11698 7984 11704
rect 7380 11688 7432 11694
rect 7380 11630 7432 11636
rect 7392 11354 7420 11630
rect 7380 11348 7432 11354
rect 7380 11290 7432 11296
rect 8404 10962 8432 12158
rect 8484 12096 8536 12102
rect 8484 12038 8536 12044
rect 8496 11082 8524 12038
rect 8576 11280 8628 11286
rect 8576 11222 8628 11228
rect 8484 11076 8536 11082
rect 8484 11018 8536 11024
rect 8404 10934 8524 10962
rect 8392 10804 8444 10810
rect 8392 10746 8444 10752
rect 7196 10736 7248 10742
rect 7196 10678 7248 10684
rect 6184 10600 6236 10606
rect 6184 10542 6236 10548
rect 6736 10600 6788 10606
rect 6736 10542 6788 10548
rect 7208 9722 7236 10678
rect 8404 10062 8432 10746
rect 8496 10588 8524 10934
rect 8588 10810 8616 11222
rect 8680 10810 8708 12174
rect 8944 11688 8996 11694
rect 8944 11630 8996 11636
rect 8956 10962 8984 11630
rect 9048 11150 9076 12854
rect 9692 12782 9720 15966
rect 9772 12980 9824 12986
rect 9772 12922 9824 12928
rect 9680 12776 9732 12782
rect 9680 12718 9732 12724
rect 9680 12368 9732 12374
rect 9680 12310 9732 12316
rect 9036 11144 9088 11150
rect 9036 11086 9088 11092
rect 8956 10934 9076 10962
rect 8576 10804 8628 10810
rect 8576 10746 8628 10752
rect 8668 10804 8720 10810
rect 8668 10746 8720 10752
rect 8576 10600 8628 10606
rect 8496 10560 8576 10588
rect 8496 10266 8524 10560
rect 8576 10542 8628 10548
rect 9048 10538 9076 10934
rect 9036 10532 9088 10538
rect 9036 10474 9088 10480
rect 8760 10464 8812 10470
rect 8760 10406 8812 10412
rect 8852 10464 8904 10470
rect 8852 10406 8904 10412
rect 8484 10260 8536 10266
rect 8484 10202 8536 10208
rect 8392 10056 8444 10062
rect 8392 9998 8444 10004
rect 7932 9920 7984 9926
rect 7932 9862 7984 9868
rect 7196 9716 7248 9722
rect 7196 9658 7248 9664
rect 7288 9580 7340 9586
rect 7288 9522 7340 9528
rect 6920 9512 6972 9518
rect 6920 9454 6972 9460
rect 6000 8492 6052 8498
rect 6000 8434 6052 8440
rect 6012 7546 6040 8434
rect 6644 8424 6696 8430
rect 6644 8366 6696 8372
rect 6552 8288 6604 8294
rect 6552 8230 6604 8236
rect 6564 7546 6592 8230
rect 6000 7540 6052 7546
rect 6000 7482 6052 7488
rect 6552 7540 6604 7546
rect 6552 7482 6604 7488
rect 5908 7472 5960 7478
rect 5908 7414 5960 7420
rect 5816 6724 5868 6730
rect 5816 6666 5868 6672
rect 5908 6724 5960 6730
rect 5908 6666 5960 6672
rect 5920 6458 5948 6666
rect 6656 6662 6684 8366
rect 6736 7744 6788 7750
rect 6736 7686 6788 7692
rect 6748 7410 6776 7686
rect 6932 7478 6960 9454
rect 7300 9178 7328 9522
rect 7288 9172 7340 9178
rect 7288 9114 7340 9120
rect 7944 8974 7972 9862
rect 8404 9722 8432 9998
rect 8576 9920 8628 9926
rect 8576 9862 8628 9868
rect 8392 9716 8444 9722
rect 8392 9658 8444 9664
rect 7932 8968 7984 8974
rect 7932 8910 7984 8916
rect 8588 8838 8616 9862
rect 8772 9110 8800 10406
rect 8864 10266 8892 10406
rect 8852 10260 8904 10266
rect 8852 10202 8904 10208
rect 9048 9674 9076 10474
rect 8864 9646 9076 9674
rect 8760 9104 8812 9110
rect 8760 9046 8812 9052
rect 8576 8832 8628 8838
rect 8576 8774 8628 8780
rect 8392 8492 8444 8498
rect 8392 8434 8444 8440
rect 8300 8356 8352 8362
rect 8300 8298 8352 8304
rect 7288 7880 7340 7886
rect 7288 7822 7340 7828
rect 6920 7472 6972 7478
rect 6920 7414 6972 7420
rect 6736 7404 6788 7410
rect 6736 7346 6788 7352
rect 6932 6798 6960 7414
rect 7300 7342 7328 7822
rect 7472 7744 7524 7750
rect 7472 7686 7524 7692
rect 7288 7336 7340 7342
rect 7288 7278 7340 7284
rect 7196 7200 7248 7206
rect 7196 7142 7248 7148
rect 6920 6792 6972 6798
rect 6920 6734 6972 6740
rect 6644 6656 6696 6662
rect 6644 6598 6696 6604
rect 5908 6452 5960 6458
rect 5908 6394 5960 6400
rect 5448 6316 5500 6322
rect 5448 6258 5500 6264
rect 5724 6316 5776 6322
rect 5724 6258 5776 6264
rect 5736 5914 5764 6258
rect 5724 5908 5776 5914
rect 5724 5850 5776 5856
rect 5356 5636 5408 5642
rect 5356 5578 5408 5584
rect 4920 5468 5296 5477
rect 4976 5466 5000 5468
rect 5056 5466 5080 5468
rect 5136 5466 5160 5468
rect 5216 5466 5240 5468
rect 4976 5414 4986 5466
rect 5230 5414 5240 5466
rect 4976 5412 5000 5414
rect 5056 5412 5080 5414
rect 5136 5412 5160 5414
rect 5216 5412 5240 5414
rect 4920 5403 5296 5412
rect 4180 4924 4556 4933
rect 4236 4922 4260 4924
rect 4316 4922 4340 4924
rect 4396 4922 4420 4924
rect 4476 4922 4500 4924
rect 4236 4870 4246 4922
rect 4490 4870 4500 4922
rect 4236 4868 4260 4870
rect 4316 4868 4340 4870
rect 4396 4868 4420 4870
rect 4476 4868 4500 4870
rect 4180 4859 4556 4868
rect 6932 4690 6960 6734
rect 7208 6458 7236 7142
rect 7196 6452 7248 6458
rect 7196 6394 7248 6400
rect 7484 6186 7512 7686
rect 7748 7336 7800 7342
rect 7748 7278 7800 7284
rect 8208 7336 8260 7342
rect 8208 7278 8260 7284
rect 7472 6180 7524 6186
rect 7472 6122 7524 6128
rect 7484 5642 7512 6122
rect 7760 5778 7788 7278
rect 8220 6934 8248 7278
rect 8208 6928 8260 6934
rect 8208 6870 8260 6876
rect 8312 6662 8340 8298
rect 8300 6656 8352 6662
rect 8300 6598 8352 6604
rect 8312 6322 8340 6598
rect 8300 6316 8352 6322
rect 8300 6258 8352 6264
rect 7840 6112 7892 6118
rect 7840 6054 7892 6060
rect 7852 5914 7880 6054
rect 7840 5908 7892 5914
rect 7840 5850 7892 5856
rect 7748 5772 7800 5778
rect 7748 5714 7800 5720
rect 7472 5636 7524 5642
rect 7472 5578 7524 5584
rect 8024 5228 8076 5234
rect 8024 5170 8076 5176
rect 7288 5024 7340 5030
rect 7288 4966 7340 4972
rect 6920 4684 6972 4690
rect 6920 4626 6972 4632
rect 4920 4380 5296 4389
rect 4976 4378 5000 4380
rect 5056 4378 5080 4380
rect 5136 4378 5160 4380
rect 5216 4378 5240 4380
rect 4976 4326 4986 4378
rect 5230 4326 5240 4378
rect 4976 4324 5000 4326
rect 5056 4324 5080 4326
rect 5136 4324 5160 4326
rect 5216 4324 5240 4326
rect 4920 4315 5296 4324
rect 6932 4146 6960 4626
rect 7300 4622 7328 4966
rect 8036 4826 8064 5170
rect 8024 4820 8076 4826
rect 8024 4762 8076 4768
rect 8404 4690 8432 8434
rect 8484 8356 8536 8362
rect 8484 8298 8536 8304
rect 8496 6254 8524 8298
rect 8588 7698 8616 8774
rect 8668 8288 8720 8294
rect 8668 8230 8720 8236
rect 8680 7886 8708 8230
rect 8668 7880 8720 7886
rect 8668 7822 8720 7828
rect 8588 7670 8708 7698
rect 8576 7336 8628 7342
rect 8576 7278 8628 7284
rect 8588 6322 8616 7278
rect 8576 6316 8628 6322
rect 8576 6258 8628 6264
rect 8484 6248 8536 6254
rect 8484 6190 8536 6196
rect 8680 5370 8708 7670
rect 8864 7478 8892 9646
rect 9692 8650 9720 12310
rect 9784 12238 9812 12922
rect 9968 12306 9996 18550
rect 10180 17980 10556 17989
rect 10236 17978 10260 17980
rect 10316 17978 10340 17980
rect 10396 17978 10420 17980
rect 10476 17978 10500 17980
rect 10236 17926 10246 17978
rect 10490 17926 10500 17978
rect 10236 17924 10260 17926
rect 10316 17924 10340 17926
rect 10396 17924 10420 17926
rect 10476 17924 10500 17926
rect 10180 17915 10556 17924
rect 10600 17196 10652 17202
rect 10600 17138 10652 17144
rect 10048 16992 10100 16998
rect 10048 16934 10100 16940
rect 10060 16590 10088 16934
rect 10180 16892 10556 16901
rect 10236 16890 10260 16892
rect 10316 16890 10340 16892
rect 10396 16890 10420 16892
rect 10476 16890 10500 16892
rect 10236 16838 10246 16890
rect 10490 16838 10500 16890
rect 10236 16836 10260 16838
rect 10316 16836 10340 16838
rect 10396 16836 10420 16838
rect 10476 16836 10500 16838
rect 10180 16827 10556 16836
rect 10048 16584 10100 16590
rect 10048 16526 10100 16532
rect 10612 16250 10640 17138
rect 10600 16244 10652 16250
rect 10600 16186 10652 16192
rect 10692 16040 10744 16046
rect 10692 15982 10744 15988
rect 10600 15904 10652 15910
rect 10600 15846 10652 15852
rect 10180 15804 10556 15813
rect 10236 15802 10260 15804
rect 10316 15802 10340 15804
rect 10396 15802 10420 15804
rect 10476 15802 10500 15804
rect 10236 15750 10246 15802
rect 10490 15750 10500 15802
rect 10236 15748 10260 15750
rect 10316 15748 10340 15750
rect 10396 15748 10420 15750
rect 10476 15748 10500 15750
rect 10180 15739 10556 15748
rect 10416 15496 10468 15502
rect 10416 15438 10468 15444
rect 10428 15162 10456 15438
rect 10416 15156 10468 15162
rect 10416 15098 10468 15104
rect 10180 14716 10556 14725
rect 10236 14714 10260 14716
rect 10316 14714 10340 14716
rect 10396 14714 10420 14716
rect 10476 14714 10500 14716
rect 10236 14662 10246 14714
rect 10490 14662 10500 14714
rect 10236 14660 10260 14662
rect 10316 14660 10340 14662
rect 10396 14660 10420 14662
rect 10476 14660 10500 14662
rect 10180 14651 10556 14660
rect 10180 13628 10556 13637
rect 10236 13626 10260 13628
rect 10316 13626 10340 13628
rect 10396 13626 10420 13628
rect 10476 13626 10500 13628
rect 10236 13574 10246 13626
rect 10490 13574 10500 13626
rect 10236 13572 10260 13574
rect 10316 13572 10340 13574
rect 10396 13572 10420 13574
rect 10476 13572 10500 13574
rect 10180 13563 10556 13572
rect 10048 12708 10100 12714
rect 10048 12650 10100 12656
rect 10060 12374 10088 12650
rect 10180 12540 10556 12549
rect 10236 12538 10260 12540
rect 10316 12538 10340 12540
rect 10396 12538 10420 12540
rect 10476 12538 10500 12540
rect 10236 12486 10246 12538
rect 10490 12486 10500 12538
rect 10236 12484 10260 12486
rect 10316 12484 10340 12486
rect 10396 12484 10420 12486
rect 10476 12484 10500 12486
rect 10180 12475 10556 12484
rect 10048 12368 10100 12374
rect 10048 12310 10100 12316
rect 9956 12300 10008 12306
rect 9956 12242 10008 12248
rect 9772 12232 9824 12238
rect 9772 12174 9824 12180
rect 9968 11914 9996 12242
rect 10048 12096 10100 12102
rect 10048 12038 10100 12044
rect 9784 11886 9996 11914
rect 9784 10146 9812 11886
rect 9864 11756 9916 11762
rect 9864 11698 9916 11704
rect 9876 11082 9904 11698
rect 9864 11076 9916 11082
rect 9864 11018 9916 11024
rect 9956 11008 10008 11014
rect 9956 10950 10008 10956
rect 9968 10810 9996 10950
rect 9956 10804 10008 10810
rect 9956 10746 10008 10752
rect 10060 10266 10088 12038
rect 10180 11452 10556 11461
rect 10236 11450 10260 11452
rect 10316 11450 10340 11452
rect 10396 11450 10420 11452
rect 10476 11450 10500 11452
rect 10236 11398 10246 11450
rect 10490 11398 10500 11450
rect 10236 11396 10260 11398
rect 10316 11396 10340 11398
rect 10396 11396 10420 11398
rect 10476 11396 10500 11398
rect 10180 11387 10556 11396
rect 10180 10364 10556 10373
rect 10236 10362 10260 10364
rect 10316 10362 10340 10364
rect 10396 10362 10420 10364
rect 10476 10362 10500 10364
rect 10236 10310 10246 10362
rect 10490 10310 10500 10362
rect 10236 10308 10260 10310
rect 10316 10308 10340 10310
rect 10396 10308 10420 10310
rect 10476 10308 10500 10310
rect 10180 10299 10556 10308
rect 10048 10260 10100 10266
rect 10048 10202 10100 10208
rect 9784 10118 10088 10146
rect 9864 9988 9916 9994
rect 9864 9930 9916 9936
rect 9772 8968 9824 8974
rect 9772 8910 9824 8916
rect 9416 8622 9720 8650
rect 8944 8492 8996 8498
rect 8944 8434 8996 8440
rect 9220 8492 9272 8498
rect 9220 8434 9272 8440
rect 8852 7472 8904 7478
rect 8852 7414 8904 7420
rect 8760 7404 8812 7410
rect 8760 7346 8812 7352
rect 8772 7002 8800 7346
rect 8760 6996 8812 7002
rect 8760 6938 8812 6944
rect 8956 6322 8984 8434
rect 9232 6458 9260 8434
rect 9312 8356 9364 8362
rect 9312 8298 9364 8304
rect 9324 7886 9352 8298
rect 9312 7880 9364 7886
rect 9312 7822 9364 7828
rect 9416 7290 9444 8622
rect 9680 8492 9732 8498
rect 9680 8434 9732 8440
rect 9692 7886 9720 8434
rect 9784 8090 9812 8910
rect 9876 8634 9904 9930
rect 9864 8628 9916 8634
rect 9864 8570 9916 8576
rect 9956 8560 10008 8566
rect 10060 8537 10088 10118
rect 10180 9276 10556 9285
rect 10236 9274 10260 9276
rect 10316 9274 10340 9276
rect 10396 9274 10420 9276
rect 10476 9274 10500 9276
rect 10236 9222 10246 9274
rect 10490 9222 10500 9274
rect 10236 9220 10260 9222
rect 10316 9220 10340 9222
rect 10396 9220 10420 9222
rect 10476 9220 10500 9222
rect 10180 9211 10556 9220
rect 10324 8832 10376 8838
rect 10324 8774 10376 8780
rect 9956 8502 10008 8508
rect 10046 8528 10102 8537
rect 9864 8288 9916 8294
rect 9864 8230 9916 8236
rect 9772 8084 9824 8090
rect 9772 8026 9824 8032
rect 9876 7970 9904 8230
rect 9784 7942 9904 7970
rect 9680 7880 9732 7886
rect 9680 7822 9732 7828
rect 9784 7818 9812 7942
rect 9772 7812 9824 7818
rect 9772 7754 9824 7760
rect 9680 7472 9732 7478
rect 9678 7440 9680 7449
rect 9732 7440 9734 7449
rect 9678 7375 9734 7384
rect 9416 7262 9720 7290
rect 9588 6792 9640 6798
rect 9588 6734 9640 6740
rect 9220 6452 9272 6458
rect 9220 6394 9272 6400
rect 9600 6322 9628 6734
rect 8852 6316 8904 6322
rect 8852 6258 8904 6264
rect 8944 6316 8996 6322
rect 8944 6258 8996 6264
rect 9588 6316 9640 6322
rect 9588 6258 9640 6264
rect 8668 5364 8720 5370
rect 8668 5306 8720 5312
rect 8864 5098 8892 6258
rect 8852 5092 8904 5098
rect 8852 5034 8904 5040
rect 8864 4758 8892 5034
rect 9220 5024 9272 5030
rect 9220 4966 9272 4972
rect 9232 4826 9260 4966
rect 9220 4820 9272 4826
rect 9220 4762 9272 4768
rect 8852 4752 8904 4758
rect 8852 4694 8904 4700
rect 8392 4684 8444 4690
rect 8392 4626 8444 4632
rect 7288 4616 7340 4622
rect 7288 4558 7340 4564
rect 7288 4480 7340 4486
rect 7288 4422 7340 4428
rect 7300 4282 7328 4422
rect 8404 4282 8432 4626
rect 7288 4276 7340 4282
rect 7288 4218 7340 4224
rect 8392 4276 8444 4282
rect 8392 4218 8444 4224
rect 6920 4140 6972 4146
rect 6920 4082 6972 4088
rect 4180 3836 4556 3845
rect 4236 3834 4260 3836
rect 4316 3834 4340 3836
rect 4396 3834 4420 3836
rect 4476 3834 4500 3836
rect 4236 3782 4246 3834
rect 4490 3782 4500 3834
rect 4236 3780 4260 3782
rect 4316 3780 4340 3782
rect 4396 3780 4420 3782
rect 4476 3780 4500 3782
rect 4180 3771 4556 3780
rect 4920 3292 5296 3301
rect 4976 3290 5000 3292
rect 5056 3290 5080 3292
rect 5136 3290 5160 3292
rect 5216 3290 5240 3292
rect 4976 3238 4986 3290
rect 5230 3238 5240 3290
rect 4976 3236 5000 3238
rect 5056 3236 5080 3238
rect 5136 3236 5160 3238
rect 5216 3236 5240 3238
rect 4920 3227 5296 3236
rect 6932 3058 6960 4082
rect 9692 4026 9720 7262
rect 9784 6866 9812 7754
rect 9968 7546 9996 8502
rect 10046 8463 10102 8472
rect 10336 8430 10364 8774
rect 10324 8424 10376 8430
rect 10324 8366 10376 8372
rect 10048 8356 10100 8362
rect 10048 8298 10100 8304
rect 9956 7540 10008 7546
rect 10060 7528 10088 8298
rect 10180 8188 10556 8197
rect 10236 8186 10260 8188
rect 10316 8186 10340 8188
rect 10396 8186 10420 8188
rect 10476 8186 10500 8188
rect 10236 8134 10246 8186
rect 10490 8134 10500 8186
rect 10236 8132 10260 8134
rect 10316 8132 10340 8134
rect 10396 8132 10420 8134
rect 10476 8132 10500 8134
rect 10180 8123 10556 8132
rect 10508 7812 10560 7818
rect 10508 7754 10560 7760
rect 10520 7546 10548 7754
rect 10508 7540 10560 7546
rect 10060 7500 10180 7528
rect 9956 7482 10008 7488
rect 10152 7188 10180 7500
rect 10508 7482 10560 7488
rect 10060 7160 10180 7188
rect 9772 6860 9824 6866
rect 9772 6802 9824 6808
rect 9770 6760 9826 6769
rect 10060 6730 10088 7160
rect 10180 7100 10556 7109
rect 10236 7098 10260 7100
rect 10316 7098 10340 7100
rect 10396 7098 10420 7100
rect 10476 7098 10500 7100
rect 10236 7046 10246 7098
rect 10490 7046 10500 7098
rect 10236 7044 10260 7046
rect 10316 7044 10340 7046
rect 10396 7044 10420 7046
rect 10476 7044 10500 7046
rect 10180 7035 10556 7044
rect 9770 6695 9826 6704
rect 10048 6724 10100 6730
rect 9784 6662 9812 6695
rect 10048 6666 10100 6672
rect 9772 6656 9824 6662
rect 9772 6598 9824 6604
rect 9784 5370 9812 6598
rect 10180 6012 10556 6021
rect 10236 6010 10260 6012
rect 10316 6010 10340 6012
rect 10396 6010 10420 6012
rect 10476 6010 10500 6012
rect 10236 5958 10246 6010
rect 10490 5958 10500 6010
rect 10236 5956 10260 5958
rect 10316 5956 10340 5958
rect 10396 5956 10420 5958
rect 10476 5956 10500 5958
rect 10180 5947 10556 5956
rect 9772 5364 9824 5370
rect 9772 5306 9824 5312
rect 10046 4992 10102 5001
rect 10046 4927 10102 4936
rect 10060 4078 10088 4927
rect 10180 4924 10556 4933
rect 10236 4922 10260 4924
rect 10316 4922 10340 4924
rect 10396 4922 10420 4924
rect 10476 4922 10500 4924
rect 10236 4870 10246 4922
rect 10490 4870 10500 4922
rect 10236 4868 10260 4870
rect 10316 4868 10340 4870
rect 10396 4868 10420 4870
rect 10476 4868 10500 4870
rect 10180 4859 10556 4868
rect 10508 4480 10560 4486
rect 10508 4422 10560 4428
rect 10520 4282 10548 4422
rect 10508 4276 10560 4282
rect 10508 4218 10560 4224
rect 10612 4146 10640 15846
rect 10704 15094 10732 15982
rect 10796 15978 10824 20538
rect 11520 20392 11572 20398
rect 11520 20334 11572 20340
rect 11336 19712 11388 19718
rect 11336 19654 11388 19660
rect 10920 19612 11296 19621
rect 10976 19610 11000 19612
rect 11056 19610 11080 19612
rect 11136 19610 11160 19612
rect 11216 19610 11240 19612
rect 10976 19558 10986 19610
rect 11230 19558 11240 19610
rect 10976 19556 11000 19558
rect 11056 19556 11080 19558
rect 11136 19556 11160 19558
rect 11216 19556 11240 19558
rect 10920 19547 11296 19556
rect 11348 18766 11376 19654
rect 11532 19378 11560 20334
rect 11520 19372 11572 19378
rect 11520 19314 11572 19320
rect 11532 18834 11560 19314
rect 11624 18970 11652 25706
rect 12164 25696 12216 25702
rect 12164 25638 12216 25644
rect 12072 25356 12124 25362
rect 12072 25298 12124 25304
rect 12084 24138 12112 25298
rect 12176 24750 12204 25638
rect 12256 25152 12308 25158
rect 12256 25094 12308 25100
rect 12268 24954 12296 25094
rect 12256 24948 12308 24954
rect 12256 24890 12308 24896
rect 12164 24744 12216 24750
rect 12216 24704 12296 24732
rect 12164 24686 12216 24692
rect 12164 24608 12216 24614
rect 12164 24550 12216 24556
rect 12176 24410 12204 24550
rect 12164 24404 12216 24410
rect 12164 24346 12216 24352
rect 12072 24132 12124 24138
rect 12072 24074 12124 24080
rect 12164 24132 12216 24138
rect 12164 24074 12216 24080
rect 12176 22438 12204 24074
rect 12164 22432 12216 22438
rect 12164 22374 12216 22380
rect 12268 21010 12296 24704
rect 12348 24404 12400 24410
rect 12348 24346 12400 24352
rect 12360 23662 12388 24346
rect 12544 23866 12572 26862
rect 12808 26852 12860 26858
rect 12808 26794 12860 26800
rect 12716 24064 12768 24070
rect 12716 24006 12768 24012
rect 12532 23860 12584 23866
rect 12532 23802 12584 23808
rect 12348 23656 12400 23662
rect 12348 23598 12400 23604
rect 12728 21690 12756 24006
rect 12820 22982 12848 26794
rect 12992 24200 13044 24206
rect 12992 24142 13044 24148
rect 13004 23662 13032 24142
rect 12992 23656 13044 23662
rect 12992 23598 13044 23604
rect 13004 23050 13032 23598
rect 12992 23044 13044 23050
rect 12992 22986 13044 22992
rect 12808 22976 12860 22982
rect 12808 22918 12860 22924
rect 12716 21684 12768 21690
rect 12716 21626 12768 21632
rect 12820 21418 12848 22918
rect 13004 22574 13032 22986
rect 12992 22568 13044 22574
rect 12992 22510 13044 22516
rect 12808 21412 12860 21418
rect 12808 21354 12860 21360
rect 12532 21140 12584 21146
rect 12532 21082 12584 21088
rect 12256 21004 12308 21010
rect 12256 20946 12308 20952
rect 12164 20936 12216 20942
rect 12164 20878 12216 20884
rect 12176 20777 12204 20878
rect 12162 20768 12218 20777
rect 12162 20703 12218 20712
rect 12544 20330 12572 21082
rect 12900 20868 12952 20874
rect 12900 20810 12952 20816
rect 12624 20800 12676 20806
rect 12624 20742 12676 20748
rect 12532 20324 12584 20330
rect 12532 20266 12584 20272
rect 12348 20256 12400 20262
rect 12348 20198 12400 20204
rect 12164 19848 12216 19854
rect 12164 19790 12216 19796
rect 12256 19848 12308 19854
rect 12256 19790 12308 19796
rect 12072 19712 12124 19718
rect 12072 19654 12124 19660
rect 12084 19514 12112 19654
rect 12072 19508 12124 19514
rect 12072 19450 12124 19456
rect 12176 19378 12204 19790
rect 12164 19372 12216 19378
rect 12164 19314 12216 19320
rect 11612 18964 11664 18970
rect 11612 18906 11664 18912
rect 11980 18964 12032 18970
rect 11980 18906 12032 18912
rect 11520 18828 11572 18834
rect 11520 18770 11572 18776
rect 11336 18760 11388 18766
rect 11336 18702 11388 18708
rect 11888 18692 11940 18698
rect 11888 18634 11940 18640
rect 10920 18524 11296 18533
rect 10976 18522 11000 18524
rect 11056 18522 11080 18524
rect 11136 18522 11160 18524
rect 11216 18522 11240 18524
rect 10976 18470 10986 18522
rect 11230 18470 11240 18522
rect 10976 18468 11000 18470
rect 11056 18468 11080 18470
rect 11136 18468 11160 18470
rect 11216 18468 11240 18470
rect 10920 18459 11296 18468
rect 11900 18426 11928 18634
rect 11888 18420 11940 18426
rect 11888 18362 11940 18368
rect 10920 17436 11296 17445
rect 10976 17434 11000 17436
rect 11056 17434 11080 17436
rect 11136 17434 11160 17436
rect 11216 17434 11240 17436
rect 10976 17382 10986 17434
rect 11230 17382 11240 17434
rect 10976 17380 11000 17382
rect 11056 17380 11080 17382
rect 11136 17380 11160 17382
rect 11216 17380 11240 17382
rect 10920 17371 11296 17380
rect 11704 16720 11756 16726
rect 11704 16662 11756 16668
rect 11992 16674 12020 18906
rect 12176 17678 12204 19314
rect 12268 18426 12296 19790
rect 12256 18420 12308 18426
rect 12256 18362 12308 18368
rect 12164 17672 12216 17678
rect 12164 17614 12216 17620
rect 12360 17610 12388 20198
rect 12440 19440 12492 19446
rect 12440 19382 12492 19388
rect 12452 17678 12480 19382
rect 12544 17678 12572 20266
rect 12636 17746 12664 20742
rect 12912 20398 12940 20810
rect 12900 20392 12952 20398
rect 12900 20334 12952 20340
rect 12900 19848 12952 19854
rect 12900 19790 12952 19796
rect 12808 19712 12860 19718
rect 12808 19654 12860 19660
rect 12820 18426 12848 19654
rect 12912 19514 12940 19790
rect 12900 19508 12952 19514
rect 12900 19450 12952 19456
rect 12992 19168 13044 19174
rect 12992 19110 13044 19116
rect 12808 18420 12860 18426
rect 12808 18362 12860 18368
rect 12900 18420 12952 18426
rect 12900 18362 12952 18368
rect 12912 18222 12940 18362
rect 13004 18290 13032 19110
rect 12992 18284 13044 18290
rect 12992 18226 13044 18232
rect 12900 18216 12952 18222
rect 12900 18158 12952 18164
rect 12624 17740 12676 17746
rect 12624 17682 12676 17688
rect 12440 17672 12492 17678
rect 12440 17614 12492 17620
rect 12532 17672 12584 17678
rect 12532 17614 12584 17620
rect 12348 17604 12400 17610
rect 12348 17546 12400 17552
rect 12072 16992 12124 16998
rect 12072 16934 12124 16940
rect 12084 16794 12112 16934
rect 12072 16788 12124 16794
rect 12072 16730 12124 16736
rect 11336 16448 11388 16454
rect 11336 16390 11388 16396
rect 10920 16348 11296 16357
rect 10976 16346 11000 16348
rect 11056 16346 11080 16348
rect 11136 16346 11160 16348
rect 11216 16346 11240 16348
rect 10976 16294 10986 16346
rect 11230 16294 11240 16346
rect 10976 16292 11000 16294
rect 11056 16292 11080 16294
rect 11136 16292 11160 16294
rect 11216 16292 11240 16294
rect 10920 16283 11296 16292
rect 11348 16250 11376 16390
rect 11336 16244 11388 16250
rect 11336 16186 11388 16192
rect 11716 16182 11744 16662
rect 11992 16646 12112 16674
rect 11704 16176 11756 16182
rect 11704 16118 11756 16124
rect 11796 16108 11848 16114
rect 11796 16050 11848 16056
rect 10784 15972 10836 15978
rect 10784 15914 10836 15920
rect 10920 15260 11296 15269
rect 10976 15258 11000 15260
rect 11056 15258 11080 15260
rect 11136 15258 11160 15260
rect 11216 15258 11240 15260
rect 10976 15206 10986 15258
rect 11230 15206 11240 15258
rect 10976 15204 11000 15206
rect 11056 15204 11080 15206
rect 11136 15204 11160 15206
rect 11216 15204 11240 15206
rect 10920 15195 11296 15204
rect 10692 15088 10744 15094
rect 10692 15030 10744 15036
rect 10784 14272 10836 14278
rect 10784 14214 10836 14220
rect 10796 14074 10824 14214
rect 10920 14172 11296 14181
rect 10976 14170 11000 14172
rect 11056 14170 11080 14172
rect 11136 14170 11160 14172
rect 11216 14170 11240 14172
rect 10976 14118 10986 14170
rect 11230 14118 11240 14170
rect 10976 14116 11000 14118
rect 11056 14116 11080 14118
rect 11136 14116 11160 14118
rect 11216 14116 11240 14118
rect 10920 14107 11296 14116
rect 10784 14068 10836 14074
rect 10784 14010 10836 14016
rect 10920 13084 11296 13093
rect 10976 13082 11000 13084
rect 11056 13082 11080 13084
rect 11136 13082 11160 13084
rect 11216 13082 11240 13084
rect 10976 13030 10986 13082
rect 11230 13030 11240 13082
rect 10976 13028 11000 13030
rect 11056 13028 11080 13030
rect 11136 13028 11160 13030
rect 11216 13028 11240 13030
rect 10920 13019 11296 13028
rect 10920 11996 11296 12005
rect 10976 11994 11000 11996
rect 11056 11994 11080 11996
rect 11136 11994 11160 11996
rect 11216 11994 11240 11996
rect 10976 11942 10986 11994
rect 11230 11942 11240 11994
rect 10976 11940 11000 11942
rect 11056 11940 11080 11942
rect 11136 11940 11160 11942
rect 11216 11940 11240 11942
rect 10920 11931 11296 11940
rect 11336 11212 11388 11218
rect 11336 11154 11388 11160
rect 10692 11008 10744 11014
rect 10692 10950 10744 10956
rect 10704 10742 10732 10950
rect 10920 10908 11296 10917
rect 10976 10906 11000 10908
rect 11056 10906 11080 10908
rect 11136 10906 11160 10908
rect 11216 10906 11240 10908
rect 10976 10854 10986 10906
rect 11230 10854 11240 10906
rect 10976 10852 11000 10854
rect 11056 10852 11080 10854
rect 11136 10852 11160 10854
rect 11216 10852 11240 10854
rect 10920 10843 11296 10852
rect 11348 10810 11376 11154
rect 11520 11144 11572 11150
rect 11520 11086 11572 11092
rect 11532 10810 11560 11086
rect 11336 10804 11388 10810
rect 11336 10746 11388 10752
rect 11520 10804 11572 10810
rect 11520 10746 11572 10752
rect 10692 10736 10744 10742
rect 10692 10678 10744 10684
rect 10876 10736 10928 10742
rect 10876 10678 10928 10684
rect 10888 10010 10916 10678
rect 11348 10062 11376 10746
rect 11612 10736 11664 10742
rect 11612 10678 11664 10684
rect 10796 9982 10916 10010
rect 11336 10056 11388 10062
rect 11336 9998 11388 10004
rect 10796 8945 10824 9982
rect 11520 9920 11572 9926
rect 11520 9862 11572 9868
rect 10920 9820 11296 9829
rect 10976 9818 11000 9820
rect 11056 9818 11080 9820
rect 11136 9818 11160 9820
rect 11216 9818 11240 9820
rect 10976 9766 10986 9818
rect 11230 9766 11240 9818
rect 10976 9764 11000 9766
rect 11056 9764 11080 9766
rect 11136 9764 11160 9766
rect 11216 9764 11240 9766
rect 10920 9755 11296 9764
rect 11244 9716 11296 9722
rect 11244 9658 11296 9664
rect 11152 9580 11204 9586
rect 11152 9522 11204 9528
rect 11164 9178 11192 9522
rect 11256 9194 11284 9658
rect 11152 9172 11204 9178
rect 11256 9166 11468 9194
rect 11152 9114 11204 9120
rect 11336 9104 11388 9110
rect 11336 9046 11388 9052
rect 10782 8936 10838 8945
rect 10692 8900 10744 8906
rect 10782 8871 10838 8880
rect 10692 8842 10744 8848
rect 10704 7970 10732 8842
rect 10784 8832 10836 8838
rect 10784 8774 10836 8780
rect 10796 8634 10824 8774
rect 10920 8732 11296 8741
rect 10976 8730 11000 8732
rect 11056 8730 11080 8732
rect 11136 8730 11160 8732
rect 11216 8730 11240 8732
rect 10976 8678 10986 8730
rect 11230 8678 11240 8730
rect 10976 8676 11000 8678
rect 11056 8676 11080 8678
rect 11136 8676 11160 8678
rect 11216 8676 11240 8678
rect 10920 8667 11296 8676
rect 10784 8628 10836 8634
rect 10784 8570 10836 8576
rect 10784 8424 10836 8430
rect 10784 8366 10836 8372
rect 10796 8294 10824 8366
rect 10784 8288 10836 8294
rect 10784 8230 10836 8236
rect 10704 7942 10824 7970
rect 10692 7812 10744 7818
rect 10692 7754 10744 7760
rect 10704 7002 10732 7754
rect 10692 6996 10744 7002
rect 10692 6938 10744 6944
rect 10796 4706 10824 7942
rect 11348 7886 11376 9046
rect 11336 7880 11388 7886
rect 11336 7822 11388 7828
rect 11440 7818 11468 9166
rect 11532 8974 11560 9862
rect 11624 9586 11652 10678
rect 11808 9994 11836 16050
rect 11980 15496 12032 15502
rect 11980 15438 12032 15444
rect 11888 14272 11940 14278
rect 11888 14214 11940 14220
rect 11900 13870 11928 14214
rect 11992 14074 12020 15438
rect 11980 14068 12032 14074
rect 11980 14010 12032 14016
rect 12084 13870 12112 16646
rect 12360 15366 12388 17546
rect 12544 15434 12572 17614
rect 12532 15428 12584 15434
rect 12532 15370 12584 15376
rect 12348 15360 12400 15366
rect 12348 15302 12400 15308
rect 12440 15088 12492 15094
rect 12440 15030 12492 15036
rect 12452 14618 12480 15030
rect 12544 14906 12572 15370
rect 12636 15162 12664 17682
rect 13096 16794 13124 31726
rect 13544 31690 13596 31696
rect 13556 31482 13584 31690
rect 19352 31686 19380 32370
rect 22180 32124 22556 32133
rect 22236 32122 22260 32124
rect 22316 32122 22340 32124
rect 22396 32122 22420 32124
rect 22476 32122 22500 32124
rect 22236 32070 22246 32122
rect 22490 32070 22500 32122
rect 22236 32068 22260 32070
rect 22316 32068 22340 32070
rect 22396 32068 22420 32070
rect 22476 32068 22500 32070
rect 22180 32059 22556 32068
rect 20168 31816 20220 31822
rect 20168 31758 20220 31764
rect 18236 31680 18288 31686
rect 18236 31622 18288 31628
rect 19340 31680 19392 31686
rect 19340 31622 19392 31628
rect 16920 31580 17296 31589
rect 16976 31578 17000 31580
rect 17056 31578 17080 31580
rect 17136 31578 17160 31580
rect 17216 31578 17240 31580
rect 16976 31526 16986 31578
rect 17230 31526 17240 31578
rect 16976 31524 17000 31526
rect 17056 31524 17080 31526
rect 17136 31524 17160 31526
rect 17216 31524 17240 31526
rect 16920 31515 17296 31524
rect 13544 31476 13596 31482
rect 13544 31418 13596 31424
rect 13176 31136 13228 31142
rect 13176 31078 13228 31084
rect 13188 30938 13216 31078
rect 13556 30938 13584 31418
rect 18248 31414 18276 31622
rect 14004 31408 14056 31414
rect 14004 31350 14056 31356
rect 14372 31408 14424 31414
rect 14372 31350 14424 31356
rect 14832 31408 14884 31414
rect 14832 31350 14884 31356
rect 18236 31408 18288 31414
rect 18236 31350 18288 31356
rect 19432 31408 19484 31414
rect 19432 31350 19484 31356
rect 13176 30932 13228 30938
rect 13176 30874 13228 30880
rect 13544 30932 13596 30938
rect 13544 30874 13596 30880
rect 13452 30660 13504 30666
rect 13452 30602 13504 30608
rect 13268 29504 13320 29510
rect 13268 29446 13320 29452
rect 13280 29170 13308 29446
rect 13268 29164 13320 29170
rect 13268 29106 13320 29112
rect 13464 26926 13492 30602
rect 13912 30252 13964 30258
rect 13912 30194 13964 30200
rect 13636 30048 13688 30054
rect 13636 29990 13688 29996
rect 13648 29510 13676 29990
rect 13924 29850 13952 30194
rect 14016 29850 14044 31350
rect 14096 31272 14148 31278
rect 14096 31214 14148 31220
rect 14108 30938 14136 31214
rect 14096 30932 14148 30938
rect 14096 30874 14148 30880
rect 14096 30660 14148 30666
rect 14096 30602 14148 30608
rect 14108 30054 14136 30602
rect 14384 30598 14412 31350
rect 14844 30938 14872 31350
rect 16764 31340 16816 31346
rect 16764 31282 16816 31288
rect 17224 31340 17276 31346
rect 17224 31282 17276 31288
rect 17500 31340 17552 31346
rect 17500 31282 17552 31288
rect 17868 31340 17920 31346
rect 17868 31282 17920 31288
rect 15476 31136 15528 31142
rect 15476 31078 15528 31084
rect 14832 30932 14884 30938
rect 14832 30874 14884 30880
rect 15488 30802 15516 31078
rect 16180 31036 16556 31045
rect 16236 31034 16260 31036
rect 16316 31034 16340 31036
rect 16396 31034 16420 31036
rect 16476 31034 16500 31036
rect 16236 30982 16246 31034
rect 16490 30982 16500 31034
rect 16236 30980 16260 30982
rect 16316 30980 16340 30982
rect 16396 30980 16420 30982
rect 16476 30980 16500 30982
rect 16180 30971 16556 30980
rect 15476 30796 15528 30802
rect 15476 30738 15528 30744
rect 15016 30728 15068 30734
rect 15016 30670 15068 30676
rect 14188 30592 14240 30598
rect 14188 30534 14240 30540
rect 14280 30592 14332 30598
rect 14280 30534 14332 30540
rect 14372 30592 14424 30598
rect 14372 30534 14424 30540
rect 14096 30048 14148 30054
rect 14096 29990 14148 29996
rect 13912 29844 13964 29850
rect 13912 29786 13964 29792
rect 14004 29844 14056 29850
rect 14004 29786 14056 29792
rect 13636 29504 13688 29510
rect 13636 29446 13688 29452
rect 13648 26994 13676 29446
rect 13728 29164 13780 29170
rect 13728 29106 13780 29112
rect 13740 28218 13768 29106
rect 14002 29064 14058 29073
rect 14108 29050 14136 29990
rect 14200 29646 14228 30534
rect 14292 29646 14320 30534
rect 14188 29640 14240 29646
rect 14188 29582 14240 29588
rect 14280 29640 14332 29646
rect 14280 29582 14332 29588
rect 14384 29458 14412 30534
rect 15028 30258 15056 30670
rect 15752 30660 15804 30666
rect 15752 30602 15804 30608
rect 15764 30394 15792 30602
rect 16580 30592 16632 30598
rect 16580 30534 16632 30540
rect 15752 30388 15804 30394
rect 15752 30330 15804 30336
rect 14924 30252 14976 30258
rect 14924 30194 14976 30200
rect 15016 30252 15068 30258
rect 15016 30194 15068 30200
rect 15752 30252 15804 30258
rect 15752 30194 15804 30200
rect 14648 30184 14700 30190
rect 14648 30126 14700 30132
rect 14058 29022 14136 29050
rect 14200 29430 14412 29458
rect 14002 28999 14058 29008
rect 13820 28484 13872 28490
rect 13820 28426 13872 28432
rect 13832 28218 13860 28426
rect 14004 28416 14056 28422
rect 14004 28358 14056 28364
rect 14096 28416 14148 28422
rect 14096 28358 14148 28364
rect 13728 28212 13780 28218
rect 13728 28154 13780 28160
rect 13820 28212 13872 28218
rect 13820 28154 13872 28160
rect 13912 28076 13964 28082
rect 13912 28018 13964 28024
rect 13728 28008 13780 28014
rect 13728 27950 13780 27956
rect 13636 26988 13688 26994
rect 13636 26930 13688 26936
rect 13452 26920 13504 26926
rect 13452 26862 13504 26868
rect 13176 26308 13228 26314
rect 13176 26250 13228 26256
rect 13188 25838 13216 26250
rect 13176 25832 13228 25838
rect 13176 25774 13228 25780
rect 13188 18426 13216 25774
rect 13544 24064 13596 24070
rect 13544 24006 13596 24012
rect 13636 24064 13688 24070
rect 13636 24006 13688 24012
rect 13452 23860 13504 23866
rect 13452 23802 13504 23808
rect 13464 23474 13492 23802
rect 13556 23662 13584 24006
rect 13544 23656 13596 23662
rect 13544 23598 13596 23604
rect 13648 23474 13676 24006
rect 13464 23446 13676 23474
rect 13648 23050 13676 23446
rect 13636 23044 13688 23050
rect 13636 22986 13688 22992
rect 13360 21548 13412 21554
rect 13360 21490 13412 21496
rect 13268 21344 13320 21350
rect 13268 21286 13320 21292
rect 13280 20534 13308 21286
rect 13372 20602 13400 21490
rect 13360 20596 13412 20602
rect 13360 20538 13412 20544
rect 13268 20528 13320 20534
rect 13268 20470 13320 20476
rect 13740 19310 13768 27950
rect 13924 27538 13952 28018
rect 14016 27946 14044 28358
rect 14108 28218 14136 28358
rect 14096 28212 14148 28218
rect 14096 28154 14148 28160
rect 14004 27940 14056 27946
rect 14004 27882 14056 27888
rect 14096 27872 14148 27878
rect 14096 27814 14148 27820
rect 13912 27532 13964 27538
rect 13912 27474 13964 27480
rect 14108 27470 14136 27814
rect 14096 27464 14148 27470
rect 14096 27406 14148 27412
rect 13912 26376 13964 26382
rect 13912 26318 13964 26324
rect 13924 26042 13952 26318
rect 13912 26036 13964 26042
rect 13912 25978 13964 25984
rect 13820 24744 13872 24750
rect 13872 24704 13952 24732
rect 13820 24686 13872 24692
rect 13924 24070 13952 24704
rect 14004 24676 14056 24682
rect 14004 24618 14056 24624
rect 14016 24274 14044 24618
rect 14096 24608 14148 24614
rect 14096 24550 14148 24556
rect 14004 24268 14056 24274
rect 14004 24210 14056 24216
rect 14108 24206 14136 24550
rect 14096 24200 14148 24206
rect 14096 24142 14148 24148
rect 13912 24064 13964 24070
rect 13912 24006 13964 24012
rect 13924 23730 13952 24006
rect 13912 23724 13964 23730
rect 13912 23666 13964 23672
rect 13820 23656 13872 23662
rect 14096 23656 14148 23662
rect 13872 23604 13952 23610
rect 13820 23598 13952 23604
rect 14096 23598 14148 23604
rect 13832 23582 13952 23598
rect 13924 23254 13952 23582
rect 14108 23497 14136 23598
rect 14094 23488 14150 23497
rect 14094 23423 14150 23432
rect 13912 23248 13964 23254
rect 13912 23190 13964 23196
rect 13820 23180 13872 23186
rect 13820 23122 13872 23128
rect 13832 22778 13860 23122
rect 13820 22772 13872 22778
rect 13820 22714 13872 22720
rect 13924 22642 13952 23190
rect 14096 23044 14148 23050
rect 14096 22986 14148 22992
rect 14108 22710 14136 22986
rect 14096 22704 14148 22710
rect 14096 22646 14148 22652
rect 13912 22636 13964 22642
rect 13912 22578 13964 22584
rect 14108 22574 14136 22646
rect 14096 22568 14148 22574
rect 14096 22510 14148 22516
rect 14200 20942 14228 29430
rect 14372 29164 14424 29170
rect 14372 29106 14424 29112
rect 14384 28558 14412 29106
rect 14372 28552 14424 28558
rect 14372 28494 14424 28500
rect 14384 28218 14412 28494
rect 14556 28416 14608 28422
rect 14660 28370 14688 30126
rect 14936 29850 14964 30194
rect 14924 29844 14976 29850
rect 14924 29786 14976 29792
rect 14936 28558 14964 29786
rect 15764 29510 15792 30194
rect 16180 29948 16556 29957
rect 16236 29946 16260 29948
rect 16316 29946 16340 29948
rect 16396 29946 16420 29948
rect 16476 29946 16500 29948
rect 16236 29894 16246 29946
rect 16490 29894 16500 29946
rect 16236 29892 16260 29894
rect 16316 29892 16340 29894
rect 16396 29892 16420 29894
rect 16476 29892 16500 29894
rect 16180 29883 16556 29892
rect 16028 29776 16080 29782
rect 16028 29718 16080 29724
rect 15016 29504 15068 29510
rect 15016 29446 15068 29452
rect 15752 29504 15804 29510
rect 15752 29446 15804 29452
rect 14924 28552 14976 28558
rect 14924 28494 14976 28500
rect 14740 28484 14792 28490
rect 14740 28426 14792 28432
rect 14608 28364 14688 28370
rect 14556 28358 14688 28364
rect 14568 28342 14688 28358
rect 14372 28212 14424 28218
rect 14372 28154 14424 28160
rect 14464 28212 14516 28218
rect 14464 28154 14516 28160
rect 14280 28076 14332 28082
rect 14280 28018 14332 28024
rect 14372 28076 14424 28082
rect 14476 28064 14504 28154
rect 14660 28082 14688 28342
rect 14424 28036 14504 28064
rect 14372 28018 14424 28024
rect 14292 27878 14320 28018
rect 14372 27940 14424 27946
rect 14372 27882 14424 27888
rect 14280 27872 14332 27878
rect 14280 27814 14332 27820
rect 14292 26382 14320 27814
rect 14280 26376 14332 26382
rect 14280 26318 14332 26324
rect 14384 25838 14412 27882
rect 14476 27538 14504 28036
rect 14648 28076 14700 28082
rect 14648 28018 14700 28024
rect 14464 27532 14516 27538
rect 14464 27474 14516 27480
rect 14556 27328 14608 27334
rect 14556 27270 14608 27276
rect 14568 26518 14596 27270
rect 14556 26512 14608 26518
rect 14556 26454 14608 26460
rect 14660 25906 14688 28018
rect 14752 28014 14780 28426
rect 14740 28008 14792 28014
rect 14740 27950 14792 27956
rect 14936 27674 14964 28494
rect 14924 27668 14976 27674
rect 14924 27610 14976 27616
rect 15028 27606 15056 29446
rect 15764 29102 15792 29446
rect 15752 29096 15804 29102
rect 15752 29038 15804 29044
rect 15568 27668 15620 27674
rect 15568 27610 15620 27616
rect 15016 27600 15068 27606
rect 14936 27548 15016 27554
rect 14936 27542 15068 27548
rect 14936 27526 15056 27542
rect 14832 27056 14884 27062
rect 14832 26998 14884 27004
rect 14740 26920 14792 26926
rect 14740 26862 14792 26868
rect 14752 26450 14780 26862
rect 14740 26444 14792 26450
rect 14740 26386 14792 26392
rect 14844 26042 14872 26998
rect 14936 26994 14964 27526
rect 15016 27464 15068 27470
rect 15016 27406 15068 27412
rect 15028 27130 15056 27406
rect 15016 27124 15068 27130
rect 15016 27066 15068 27072
rect 15028 26994 15056 27066
rect 14924 26988 14976 26994
rect 14924 26930 14976 26936
rect 15016 26988 15068 26994
rect 15016 26930 15068 26936
rect 15028 26874 15056 26930
rect 14936 26846 15056 26874
rect 15108 26920 15160 26926
rect 15108 26862 15160 26868
rect 14936 26518 14964 26846
rect 15016 26784 15068 26790
rect 15016 26726 15068 26732
rect 14924 26512 14976 26518
rect 14924 26454 14976 26460
rect 14936 26042 14964 26454
rect 14832 26036 14884 26042
rect 14832 25978 14884 25984
rect 14924 26036 14976 26042
rect 14924 25978 14976 25984
rect 14648 25900 14700 25906
rect 14648 25842 14700 25848
rect 14372 25832 14424 25838
rect 14372 25774 14424 25780
rect 14832 24812 14884 24818
rect 14832 24754 14884 24760
rect 14740 24200 14792 24206
rect 14740 24142 14792 24148
rect 14280 24064 14332 24070
rect 14280 24006 14332 24012
rect 14464 24064 14516 24070
rect 14464 24006 14516 24012
rect 14188 20936 14240 20942
rect 14188 20878 14240 20884
rect 14188 20800 14240 20806
rect 14188 20742 14240 20748
rect 14200 20534 14228 20742
rect 14188 20528 14240 20534
rect 14188 20470 14240 20476
rect 13452 19304 13504 19310
rect 13452 19246 13504 19252
rect 13728 19304 13780 19310
rect 13728 19246 13780 19252
rect 13268 18760 13320 18766
rect 13268 18702 13320 18708
rect 13176 18420 13228 18426
rect 13176 18362 13228 18368
rect 13280 17882 13308 18702
rect 13464 18630 13492 19246
rect 13452 18624 13504 18630
rect 13452 18566 13504 18572
rect 13268 17876 13320 17882
rect 13268 17818 13320 17824
rect 13544 17536 13596 17542
rect 13544 17478 13596 17484
rect 13556 17338 13584 17478
rect 13544 17332 13596 17338
rect 13544 17274 13596 17280
rect 13084 16788 13136 16794
rect 13084 16730 13136 16736
rect 12808 15496 12860 15502
rect 12808 15438 12860 15444
rect 12624 15156 12676 15162
rect 12624 15098 12676 15104
rect 12544 14878 12664 14906
rect 12532 14816 12584 14822
rect 12532 14758 12584 14764
rect 12440 14612 12492 14618
rect 12440 14554 12492 14560
rect 11888 13864 11940 13870
rect 11888 13806 11940 13812
rect 12072 13864 12124 13870
rect 12072 13806 12124 13812
rect 11796 9988 11848 9994
rect 11796 9930 11848 9936
rect 11612 9580 11664 9586
rect 11612 9522 11664 9528
rect 11520 8968 11572 8974
rect 11520 8910 11572 8916
rect 11624 7954 11652 9522
rect 11612 7948 11664 7954
rect 11612 7890 11664 7896
rect 11428 7812 11480 7818
rect 11428 7754 11480 7760
rect 10920 7644 11296 7653
rect 10976 7642 11000 7644
rect 11056 7642 11080 7644
rect 11136 7642 11160 7644
rect 11216 7642 11240 7644
rect 10976 7590 10986 7642
rect 11230 7590 11240 7642
rect 10976 7588 11000 7590
rect 11056 7588 11080 7590
rect 11136 7588 11160 7590
rect 11216 7588 11240 7590
rect 10920 7579 11296 7588
rect 11624 7410 11652 7890
rect 11612 7404 11664 7410
rect 11612 7346 11664 7352
rect 10876 7200 10928 7206
rect 10876 7142 10928 7148
rect 10888 6798 10916 7142
rect 10876 6792 10928 6798
rect 10876 6734 10928 6740
rect 10920 6556 11296 6565
rect 10976 6554 11000 6556
rect 11056 6554 11080 6556
rect 11136 6554 11160 6556
rect 11216 6554 11240 6556
rect 10976 6502 10986 6554
rect 11230 6502 11240 6554
rect 10976 6500 11000 6502
rect 11056 6500 11080 6502
rect 11136 6500 11160 6502
rect 11216 6500 11240 6502
rect 10920 6491 11296 6500
rect 11624 5914 11652 7346
rect 12084 7002 12112 13806
rect 12544 13326 12572 14758
rect 12532 13320 12584 13326
rect 12532 13262 12584 13268
rect 12636 12850 12664 14878
rect 12820 14278 12848 15438
rect 12900 15360 12952 15366
rect 12900 15302 12952 15308
rect 12808 14272 12860 14278
rect 12808 14214 12860 14220
rect 12820 12850 12848 14214
rect 12912 12918 12940 15302
rect 13268 15020 13320 15026
rect 13268 14962 13320 14968
rect 13280 14074 13308 14962
rect 13452 14816 13504 14822
rect 13452 14758 13504 14764
rect 13636 14816 13688 14822
rect 13636 14758 13688 14764
rect 13360 14476 13412 14482
rect 13360 14418 13412 14424
rect 13084 14068 13136 14074
rect 13084 14010 13136 14016
rect 13268 14068 13320 14074
rect 13268 14010 13320 14016
rect 12900 12912 12952 12918
rect 12900 12854 12952 12860
rect 13096 12850 13124 14010
rect 13268 12912 13320 12918
rect 13268 12854 13320 12860
rect 12624 12844 12676 12850
rect 12624 12786 12676 12792
rect 12808 12844 12860 12850
rect 12808 12786 12860 12792
rect 13084 12844 13136 12850
rect 13084 12786 13136 12792
rect 13084 11552 13136 11558
rect 13084 11494 13136 11500
rect 12990 11384 13046 11393
rect 12990 11319 13046 11328
rect 13004 11150 13032 11319
rect 12992 11144 13044 11150
rect 12992 11086 13044 11092
rect 12348 11008 12400 11014
rect 12348 10950 12400 10956
rect 12360 10810 12388 10950
rect 12348 10804 12400 10810
rect 12348 10746 12400 10752
rect 12164 10600 12216 10606
rect 12164 10542 12216 10548
rect 12176 9042 12204 10542
rect 13096 10062 13124 11494
rect 12900 10056 12952 10062
rect 12900 9998 12952 10004
rect 13084 10056 13136 10062
rect 13084 9998 13136 10004
rect 12912 9722 12940 9998
rect 12900 9716 12952 9722
rect 12900 9658 12952 9664
rect 12992 9376 13044 9382
rect 12992 9318 13044 9324
rect 12164 9036 12216 9042
rect 12164 8978 12216 8984
rect 13004 8974 13032 9318
rect 12992 8968 13044 8974
rect 12992 8910 13044 8916
rect 12440 8832 12492 8838
rect 12440 8774 12492 8780
rect 12452 8498 12480 8774
rect 12440 8492 12492 8498
rect 12440 8434 12492 8440
rect 12256 7812 12308 7818
rect 12256 7754 12308 7760
rect 12072 6996 12124 7002
rect 12072 6938 12124 6944
rect 12084 6118 12112 6938
rect 12164 6656 12216 6662
rect 12164 6598 12216 6604
rect 12176 6322 12204 6598
rect 12268 6458 12296 7754
rect 12256 6452 12308 6458
rect 12452 6440 12480 8434
rect 12532 7948 12584 7954
rect 12532 7890 12584 7896
rect 12544 7342 12572 7890
rect 12532 7336 12584 7342
rect 12532 7278 12584 7284
rect 13280 6798 13308 12854
rect 13372 8022 13400 14418
rect 13464 12918 13492 14758
rect 13648 14618 13676 14758
rect 13636 14612 13688 14618
rect 13636 14554 13688 14560
rect 13740 14498 13768 19246
rect 14292 18766 14320 24006
rect 14372 23860 14424 23866
rect 14372 23802 14424 23808
rect 14384 23118 14412 23802
rect 14372 23112 14424 23118
rect 14372 23054 14424 23060
rect 14384 22778 14412 23054
rect 14372 22772 14424 22778
rect 14372 22714 14424 22720
rect 14372 19440 14424 19446
rect 14370 19408 14372 19417
rect 14424 19408 14426 19417
rect 14370 19343 14426 19352
rect 14372 19304 14424 19310
rect 14372 19246 14424 19252
rect 14384 18970 14412 19246
rect 14372 18964 14424 18970
rect 14372 18906 14424 18912
rect 14476 18850 14504 24006
rect 14648 23792 14700 23798
rect 14648 23734 14700 23740
rect 14660 22438 14688 23734
rect 14752 23730 14780 24142
rect 14844 23798 14872 24754
rect 14832 23792 14884 23798
rect 14832 23734 14884 23740
rect 14740 23724 14792 23730
rect 14740 23666 14792 23672
rect 14752 23254 14780 23666
rect 14832 23656 14884 23662
rect 14832 23598 14884 23604
rect 14740 23248 14792 23254
rect 14740 23190 14792 23196
rect 14844 23186 14872 23598
rect 15028 23526 15056 26726
rect 15120 26450 15148 26862
rect 15384 26784 15436 26790
rect 15384 26726 15436 26732
rect 15108 26444 15160 26450
rect 15108 26386 15160 26392
rect 15200 26240 15252 26246
rect 15200 26182 15252 26188
rect 15212 25974 15240 26182
rect 15396 25974 15424 26726
rect 15580 26314 15608 27610
rect 15764 26314 15792 29038
rect 15844 27872 15896 27878
rect 15844 27814 15896 27820
rect 15856 27062 15884 27814
rect 16040 27538 16068 29718
rect 16592 29646 16620 30534
rect 16776 30410 16804 31282
rect 16856 31136 16908 31142
rect 16856 31078 16908 31084
rect 16868 30734 16896 31078
rect 17236 30818 17264 31282
rect 17316 31136 17368 31142
rect 17316 31078 17368 31084
rect 17328 30938 17356 31078
rect 17316 30932 17368 30938
rect 17316 30874 17368 30880
rect 17236 30790 17356 30818
rect 16856 30728 16908 30734
rect 16856 30670 16908 30676
rect 17328 30666 17356 30790
rect 17316 30660 17368 30666
rect 17316 30602 17368 30608
rect 16920 30492 17296 30501
rect 16976 30490 17000 30492
rect 17056 30490 17080 30492
rect 17136 30490 17160 30492
rect 17216 30490 17240 30492
rect 16976 30438 16986 30490
rect 17230 30438 17240 30490
rect 16976 30436 17000 30438
rect 17056 30436 17080 30438
rect 17136 30436 17160 30438
rect 17216 30436 17240 30438
rect 16920 30427 17296 30436
rect 16776 30382 16896 30410
rect 16672 30320 16724 30326
rect 16672 30262 16724 30268
rect 16684 29850 16712 30262
rect 16868 30054 16896 30382
rect 17328 30138 17356 30602
rect 17408 30592 17460 30598
rect 17408 30534 17460 30540
rect 17420 30258 17448 30534
rect 17512 30258 17540 31282
rect 17592 31272 17644 31278
rect 17592 31214 17644 31220
rect 17604 30938 17632 31214
rect 17776 31136 17828 31142
rect 17776 31078 17828 31084
rect 17592 30932 17644 30938
rect 17592 30874 17644 30880
rect 17592 30592 17644 30598
rect 17592 30534 17644 30540
rect 17408 30252 17460 30258
rect 17408 30194 17460 30200
rect 17500 30252 17552 30258
rect 17500 30194 17552 30200
rect 17328 30110 17448 30138
rect 16764 30048 16816 30054
rect 16764 29990 16816 29996
rect 16856 30048 16908 30054
rect 16856 29990 16908 29996
rect 16776 29850 16804 29990
rect 16672 29844 16724 29850
rect 16672 29786 16724 29792
rect 16764 29844 16816 29850
rect 16764 29786 16816 29792
rect 16580 29640 16632 29646
rect 16580 29582 16632 29588
rect 16180 28860 16556 28869
rect 16236 28858 16260 28860
rect 16316 28858 16340 28860
rect 16396 28858 16420 28860
rect 16476 28858 16500 28860
rect 16236 28806 16246 28858
rect 16490 28806 16500 28858
rect 16236 28804 16260 28806
rect 16316 28804 16340 28806
rect 16396 28804 16420 28806
rect 16476 28804 16500 28806
rect 16180 28795 16556 28804
rect 16592 28014 16620 29582
rect 16868 29510 16896 29990
rect 17420 29850 17448 30110
rect 17512 29850 17540 30194
rect 17408 29844 17460 29850
rect 17408 29786 17460 29792
rect 17500 29844 17552 29850
rect 17500 29786 17552 29792
rect 17420 29730 17448 29786
rect 17420 29714 17540 29730
rect 17420 29708 17552 29714
rect 17420 29702 17500 29708
rect 17500 29650 17552 29656
rect 17604 29578 17632 30534
rect 17788 30258 17816 31078
rect 17880 30666 17908 31282
rect 18788 31272 18840 31278
rect 18788 31214 18840 31220
rect 18512 31136 18564 31142
rect 18512 31078 18564 31084
rect 18144 30728 18196 30734
rect 18144 30670 18196 30676
rect 17868 30660 17920 30666
rect 17868 30602 17920 30608
rect 18156 30258 18184 30670
rect 18524 30258 18552 31078
rect 18800 30734 18828 31214
rect 18788 30728 18840 30734
rect 18788 30670 18840 30676
rect 19340 30728 19392 30734
rect 19340 30670 19392 30676
rect 17776 30252 17828 30258
rect 17776 30194 17828 30200
rect 18144 30252 18196 30258
rect 18144 30194 18196 30200
rect 18512 30252 18564 30258
rect 18512 30194 18564 30200
rect 17960 30048 18012 30054
rect 17960 29990 18012 29996
rect 17592 29572 17644 29578
rect 17592 29514 17644 29520
rect 16856 29504 16908 29510
rect 16856 29446 16908 29452
rect 17408 29504 17460 29510
rect 17408 29446 17460 29452
rect 16920 29404 17296 29413
rect 16976 29402 17000 29404
rect 17056 29402 17080 29404
rect 17136 29402 17160 29404
rect 17216 29402 17240 29404
rect 16976 29350 16986 29402
rect 17230 29350 17240 29402
rect 16976 29348 17000 29350
rect 17056 29348 17080 29350
rect 17136 29348 17160 29350
rect 17216 29348 17240 29350
rect 16920 29339 17296 29348
rect 16920 28316 17296 28325
rect 16976 28314 17000 28316
rect 17056 28314 17080 28316
rect 17136 28314 17160 28316
rect 17216 28314 17240 28316
rect 16976 28262 16986 28314
rect 17230 28262 17240 28314
rect 16976 28260 17000 28262
rect 17056 28260 17080 28262
rect 17136 28260 17160 28262
rect 17216 28260 17240 28262
rect 16920 28251 17296 28260
rect 16580 28008 16632 28014
rect 16948 28008 17000 28014
rect 16580 27950 16632 27956
rect 16684 27956 16948 27962
rect 16684 27950 17000 27956
rect 16684 27934 16988 27950
rect 16684 27878 16712 27934
rect 16672 27872 16724 27878
rect 16672 27814 16724 27820
rect 16764 27872 16816 27878
rect 16764 27814 16816 27820
rect 16180 27772 16556 27781
rect 16236 27770 16260 27772
rect 16316 27770 16340 27772
rect 16396 27770 16420 27772
rect 16476 27770 16500 27772
rect 16236 27718 16246 27770
rect 16490 27718 16500 27770
rect 16236 27716 16260 27718
rect 16316 27716 16340 27718
rect 16396 27716 16420 27718
rect 16476 27716 16500 27718
rect 16180 27707 16556 27716
rect 16488 27668 16540 27674
rect 16488 27610 16540 27616
rect 16028 27532 16080 27538
rect 16028 27474 16080 27480
rect 15934 27432 15990 27441
rect 15934 27367 15990 27376
rect 15948 27334 15976 27367
rect 15936 27328 15988 27334
rect 15936 27270 15988 27276
rect 15948 27062 15976 27270
rect 15844 27056 15896 27062
rect 15844 26998 15896 27004
rect 15936 27056 15988 27062
rect 15936 26998 15988 27004
rect 16040 26926 16068 27474
rect 16500 27334 16528 27610
rect 16672 27600 16724 27606
rect 16672 27542 16724 27548
rect 16120 27328 16172 27334
rect 16120 27270 16172 27276
rect 16488 27328 16540 27334
rect 16488 27270 16540 27276
rect 16580 27328 16632 27334
rect 16580 27270 16632 27276
rect 16132 26994 16160 27270
rect 16500 27112 16528 27270
rect 16408 27084 16528 27112
rect 16120 26988 16172 26994
rect 16120 26930 16172 26936
rect 16028 26920 16080 26926
rect 16132 26897 16160 26930
rect 16028 26862 16080 26868
rect 16118 26888 16174 26897
rect 16040 26450 16068 26862
rect 16408 26858 16436 27084
rect 16592 26994 16620 27270
rect 16580 26988 16632 26994
rect 16580 26930 16632 26936
rect 16118 26823 16174 26832
rect 16396 26852 16448 26858
rect 16396 26794 16448 26800
rect 16180 26684 16556 26693
rect 16236 26682 16260 26684
rect 16316 26682 16340 26684
rect 16396 26682 16420 26684
rect 16476 26682 16500 26684
rect 16236 26630 16246 26682
rect 16490 26630 16500 26682
rect 16236 26628 16260 26630
rect 16316 26628 16340 26630
rect 16396 26628 16420 26630
rect 16476 26628 16500 26630
rect 16180 26619 16556 26628
rect 16592 26466 16620 26930
rect 16028 26444 16080 26450
rect 16028 26386 16080 26392
rect 16500 26438 16620 26466
rect 15568 26308 15620 26314
rect 15568 26250 15620 26256
rect 15752 26308 15804 26314
rect 15752 26250 15804 26256
rect 16500 26246 16528 26438
rect 16488 26240 16540 26246
rect 16488 26182 16540 26188
rect 16684 26042 16712 27542
rect 16776 27402 16804 27814
rect 17420 27606 17448 29446
rect 17604 28150 17632 29514
rect 17592 28144 17644 28150
rect 17592 28086 17644 28092
rect 17684 28008 17736 28014
rect 17684 27950 17736 27956
rect 16948 27600 17000 27606
rect 16948 27542 17000 27548
rect 17408 27600 17460 27606
rect 17460 27560 17632 27588
rect 17408 27542 17460 27548
rect 16764 27396 16816 27402
rect 16764 27338 16816 27344
rect 16960 27316 16988 27542
rect 17408 27396 17460 27402
rect 17408 27338 17460 27344
rect 16868 27288 16988 27316
rect 16868 27282 16896 27288
rect 16776 27254 16896 27282
rect 16776 27062 16804 27254
rect 16920 27228 17296 27237
rect 16976 27226 17000 27228
rect 17056 27226 17080 27228
rect 17136 27226 17160 27228
rect 17216 27226 17240 27228
rect 16976 27174 16986 27226
rect 17230 27174 17240 27226
rect 16976 27172 17000 27174
rect 17056 27172 17080 27174
rect 17136 27172 17160 27174
rect 17216 27172 17240 27174
rect 16920 27163 17296 27172
rect 17040 27124 17092 27130
rect 17040 27066 17092 27072
rect 16764 27056 16816 27062
rect 16764 26998 16816 27004
rect 16776 26518 16804 26998
rect 16856 26852 16908 26858
rect 16856 26794 16908 26800
rect 16868 26761 16896 26794
rect 16854 26752 16910 26761
rect 16854 26687 16910 26696
rect 16764 26512 16816 26518
rect 16764 26454 16816 26460
rect 17052 26314 17080 27066
rect 17420 27062 17448 27338
rect 17408 27056 17460 27062
rect 17460 27016 17540 27044
rect 17408 26998 17460 27004
rect 17132 26988 17184 26994
rect 17132 26930 17184 26936
rect 17144 26897 17172 26930
rect 17130 26888 17186 26897
rect 17130 26823 17186 26832
rect 17144 26450 17172 26823
rect 17132 26444 17184 26450
rect 17132 26386 17184 26392
rect 17512 26382 17540 27016
rect 17500 26376 17552 26382
rect 17500 26318 17552 26324
rect 17604 26314 17632 27560
rect 17696 26994 17724 27950
rect 17776 27872 17828 27878
rect 17776 27814 17828 27820
rect 17788 27441 17816 27814
rect 17868 27668 17920 27674
rect 17868 27610 17920 27616
rect 17880 27470 17908 27610
rect 17868 27464 17920 27470
rect 17774 27432 17830 27441
rect 17868 27406 17920 27412
rect 17774 27367 17830 27376
rect 17788 26994 17816 27367
rect 17684 26988 17736 26994
rect 17684 26930 17736 26936
rect 17776 26988 17828 26994
rect 17776 26930 17828 26936
rect 17696 26314 17724 26930
rect 17788 26450 17816 26930
rect 17776 26444 17828 26450
rect 17776 26386 17828 26392
rect 17040 26308 17092 26314
rect 17040 26250 17092 26256
rect 17592 26308 17644 26314
rect 17592 26250 17644 26256
rect 17684 26308 17736 26314
rect 17684 26250 17736 26256
rect 16920 26140 17296 26149
rect 16976 26138 17000 26140
rect 17056 26138 17080 26140
rect 17136 26138 17160 26140
rect 17216 26138 17240 26140
rect 16976 26086 16986 26138
rect 17230 26086 17240 26138
rect 16976 26084 17000 26086
rect 17056 26084 17080 26086
rect 17136 26084 17160 26086
rect 17216 26084 17240 26086
rect 16920 26075 17296 26084
rect 16672 26036 16724 26042
rect 16672 25978 16724 25984
rect 15200 25968 15252 25974
rect 15200 25910 15252 25916
rect 15384 25968 15436 25974
rect 15384 25910 15436 25916
rect 15660 25696 15712 25702
rect 15660 25638 15712 25644
rect 15672 24410 15700 25638
rect 16180 25596 16556 25605
rect 16236 25594 16260 25596
rect 16316 25594 16340 25596
rect 16396 25594 16420 25596
rect 16476 25594 16500 25596
rect 16236 25542 16246 25594
rect 16490 25542 16500 25594
rect 16236 25540 16260 25542
rect 16316 25540 16340 25542
rect 16396 25540 16420 25542
rect 16476 25540 16500 25542
rect 16180 25531 16556 25540
rect 16488 25220 16540 25226
rect 16488 25162 16540 25168
rect 16500 24954 16528 25162
rect 16920 25052 17296 25061
rect 16976 25050 17000 25052
rect 17056 25050 17080 25052
rect 17136 25050 17160 25052
rect 17216 25050 17240 25052
rect 16976 24998 16986 25050
rect 17230 24998 17240 25050
rect 16976 24996 17000 24998
rect 17056 24996 17080 24998
rect 17136 24996 17160 24998
rect 17216 24996 17240 24998
rect 16920 24987 17296 24996
rect 16488 24948 16540 24954
rect 16488 24890 16540 24896
rect 17972 24750 18000 29990
rect 18524 29714 18552 30194
rect 18800 30190 18828 30670
rect 18788 30184 18840 30190
rect 18788 30126 18840 30132
rect 18512 29708 18564 29714
rect 18512 29650 18564 29656
rect 18052 29640 18104 29646
rect 18052 29582 18104 29588
rect 18064 28014 18092 29582
rect 18052 28008 18104 28014
rect 18052 27950 18104 27956
rect 18420 27668 18472 27674
rect 18420 27610 18472 27616
rect 18328 27600 18380 27606
rect 18328 27542 18380 27548
rect 18052 27464 18104 27470
rect 18052 27406 18104 27412
rect 18064 27130 18092 27406
rect 18340 27402 18368 27542
rect 18328 27396 18380 27402
rect 18328 27338 18380 27344
rect 18052 27124 18104 27130
rect 18052 27066 18104 27072
rect 18144 27124 18196 27130
rect 18144 27066 18196 27072
rect 18156 27010 18184 27066
rect 18064 26982 18184 27010
rect 18236 27056 18288 27062
rect 18236 26998 18288 27004
rect 18064 26897 18092 26982
rect 18050 26888 18106 26897
rect 18050 26823 18106 26832
rect 18248 26602 18276 26998
rect 18328 26988 18380 26994
rect 18328 26930 18380 26936
rect 18340 26761 18368 26930
rect 18432 26926 18460 27610
rect 18524 27470 18552 29650
rect 18880 28076 18932 28082
rect 18880 28018 18932 28024
rect 18512 27464 18564 27470
rect 18512 27406 18564 27412
rect 18420 26920 18472 26926
rect 18420 26862 18472 26868
rect 18326 26752 18382 26761
rect 18326 26687 18382 26696
rect 18156 26586 18276 26602
rect 18144 26580 18276 26586
rect 18196 26574 18276 26580
rect 18144 26522 18196 26528
rect 18236 26512 18288 26518
rect 18236 26454 18288 26460
rect 18052 26376 18104 26382
rect 18052 26318 18104 26324
rect 18064 26042 18092 26318
rect 18052 26036 18104 26042
rect 18052 25978 18104 25984
rect 18248 25906 18276 26454
rect 18328 26308 18380 26314
rect 18328 26250 18380 26256
rect 18236 25900 18288 25906
rect 18236 25842 18288 25848
rect 17960 24744 18012 24750
rect 17960 24686 18012 24692
rect 16180 24508 16556 24517
rect 16236 24506 16260 24508
rect 16316 24506 16340 24508
rect 16396 24506 16420 24508
rect 16476 24506 16500 24508
rect 16236 24454 16246 24506
rect 16490 24454 16500 24506
rect 16236 24452 16260 24454
rect 16316 24452 16340 24454
rect 16396 24452 16420 24454
rect 16476 24452 16500 24454
rect 16180 24443 16556 24452
rect 15660 24404 15712 24410
rect 15660 24346 15712 24352
rect 15292 24064 15344 24070
rect 15292 24006 15344 24012
rect 15304 23730 15332 24006
rect 15292 23724 15344 23730
rect 15292 23666 15344 23672
rect 15016 23520 15068 23526
rect 15016 23462 15068 23468
rect 15476 23520 15528 23526
rect 15476 23462 15528 23468
rect 14832 23180 14884 23186
rect 14832 23122 14884 23128
rect 15028 23118 15056 23462
rect 15488 23118 15516 23462
rect 15016 23112 15068 23118
rect 15016 23054 15068 23060
rect 15476 23112 15528 23118
rect 15476 23054 15528 23060
rect 15568 23044 15620 23050
rect 15568 22986 15620 22992
rect 15200 22976 15252 22982
rect 15200 22918 15252 22924
rect 15292 22976 15344 22982
rect 15292 22918 15344 22924
rect 15212 22438 15240 22918
rect 14648 22432 14700 22438
rect 14648 22374 14700 22380
rect 15200 22432 15252 22438
rect 15200 22374 15252 22380
rect 14924 21004 14976 21010
rect 14924 20946 14976 20952
rect 14556 20256 14608 20262
rect 14556 20198 14608 20204
rect 14384 18822 14504 18850
rect 14188 18760 14240 18766
rect 14188 18702 14240 18708
rect 14280 18760 14332 18766
rect 14280 18702 14332 18708
rect 13912 18692 13964 18698
rect 13912 18634 13964 18640
rect 13820 18624 13872 18630
rect 13820 18566 13872 18572
rect 13832 18290 13860 18566
rect 13820 18284 13872 18290
rect 13820 18226 13872 18232
rect 13556 14482 13768 14498
rect 13544 14476 13768 14482
rect 13596 14470 13768 14476
rect 13544 14418 13596 14424
rect 13728 14408 13780 14414
rect 13728 14350 13780 14356
rect 13544 14272 13596 14278
rect 13544 14214 13596 14220
rect 13556 14006 13584 14214
rect 13740 14074 13768 14350
rect 13728 14068 13780 14074
rect 13728 14010 13780 14016
rect 13544 14000 13596 14006
rect 13544 13942 13596 13948
rect 13832 12918 13860 18226
rect 13924 18086 13952 18634
rect 14200 18612 14228 18702
rect 14384 18612 14412 18822
rect 14568 18766 14596 20198
rect 14648 19440 14700 19446
rect 14648 19382 14700 19388
rect 14464 18760 14516 18766
rect 14464 18702 14516 18708
rect 14556 18760 14608 18766
rect 14556 18702 14608 18708
rect 14200 18584 14412 18612
rect 14096 18420 14148 18426
rect 14096 18362 14148 18368
rect 13912 18080 13964 18086
rect 13912 18022 13964 18028
rect 13924 17134 13952 18022
rect 14004 17536 14056 17542
rect 14004 17478 14056 17484
rect 14016 17202 14044 17478
rect 14004 17196 14056 17202
rect 14004 17138 14056 17144
rect 13912 17128 13964 17134
rect 13912 17070 13964 17076
rect 14108 17082 14136 18362
rect 14280 18284 14332 18290
rect 14280 18226 14332 18232
rect 14188 18080 14240 18086
rect 14188 18022 14240 18028
rect 14200 17202 14228 18022
rect 14292 17882 14320 18226
rect 14280 17876 14332 17882
rect 14280 17818 14332 17824
rect 14188 17196 14240 17202
rect 14188 17138 14240 17144
rect 14108 17054 14320 17082
rect 14188 16652 14240 16658
rect 14188 16594 14240 16600
rect 14096 14408 14148 14414
rect 14096 14350 14148 14356
rect 14108 13870 14136 14350
rect 14096 13864 14148 13870
rect 14096 13806 14148 13812
rect 14004 13456 14056 13462
rect 14004 13398 14056 13404
rect 14016 12986 14044 13398
rect 14108 13394 14136 13806
rect 14096 13388 14148 13394
rect 14096 13330 14148 13336
rect 14004 12980 14056 12986
rect 14004 12922 14056 12928
rect 13452 12912 13504 12918
rect 13452 12854 13504 12860
rect 13820 12912 13872 12918
rect 13820 12854 13872 12860
rect 13544 12640 13596 12646
rect 13544 12582 13596 12588
rect 13360 8016 13412 8022
rect 13360 7958 13412 7964
rect 13452 7744 13504 7750
rect 13452 7686 13504 7692
rect 13464 7410 13492 7686
rect 13452 7404 13504 7410
rect 13452 7346 13504 7352
rect 13452 7200 13504 7206
rect 13452 7142 13504 7148
rect 13464 6866 13492 7142
rect 13452 6860 13504 6866
rect 13452 6802 13504 6808
rect 13556 6798 13584 12582
rect 13728 11212 13780 11218
rect 13728 11154 13780 11160
rect 13740 11082 13768 11154
rect 13832 11098 13860 12854
rect 14108 12434 14136 13330
rect 14200 12850 14228 16594
rect 14292 13818 14320 17054
rect 14384 16658 14412 18584
rect 14476 18426 14504 18702
rect 14464 18420 14516 18426
rect 14464 18362 14516 18368
rect 14568 18222 14596 18702
rect 14556 18216 14608 18222
rect 14556 18158 14608 18164
rect 14660 16726 14688 19382
rect 14936 17746 14964 20946
rect 15016 18352 15068 18358
rect 15016 18294 15068 18300
rect 14924 17740 14976 17746
rect 14924 17682 14976 17688
rect 14648 16720 14700 16726
rect 14700 16680 14872 16708
rect 14648 16662 14700 16668
rect 14372 16652 14424 16658
rect 14372 16594 14424 16600
rect 14648 15088 14700 15094
rect 14648 15030 14700 15036
rect 14372 14816 14424 14822
rect 14372 14758 14424 14764
rect 14384 14074 14412 14758
rect 14464 14340 14516 14346
rect 14464 14282 14516 14288
rect 14476 14074 14504 14282
rect 14372 14068 14424 14074
rect 14372 14010 14424 14016
rect 14464 14068 14516 14074
rect 14464 14010 14516 14016
rect 14464 13864 14516 13870
rect 14292 13812 14464 13818
rect 14292 13806 14516 13812
rect 14292 13790 14504 13806
rect 14556 13796 14608 13802
rect 14188 12844 14240 12850
rect 14188 12786 14240 12792
rect 14016 12406 14136 12434
rect 14016 11694 14044 12406
rect 14188 11756 14240 11762
rect 14188 11698 14240 11704
rect 14004 11688 14056 11694
rect 14004 11630 14056 11636
rect 14016 11234 14044 11630
rect 14096 11552 14148 11558
rect 14096 11494 14148 11500
rect 14108 11354 14136 11494
rect 14096 11348 14148 11354
rect 14096 11290 14148 11296
rect 14016 11206 14136 11234
rect 14108 11150 14136 11206
rect 14096 11144 14148 11150
rect 13728 11076 13780 11082
rect 13832 11070 14044 11098
rect 14096 11086 14148 11092
rect 13728 11018 13780 11024
rect 13740 10588 13768 11018
rect 13820 11008 13872 11014
rect 13820 10950 13872 10956
rect 13832 10742 13860 10950
rect 13820 10736 13872 10742
rect 13820 10678 13872 10684
rect 13740 10560 13860 10588
rect 13832 9586 13860 10560
rect 13820 9580 13872 9586
rect 13820 9522 13872 9528
rect 13820 8832 13872 8838
rect 13820 8774 13872 8780
rect 13832 8634 13860 8774
rect 14016 8634 14044 11070
rect 14200 10810 14228 11698
rect 14188 10804 14240 10810
rect 14188 10746 14240 10752
rect 14096 10464 14148 10470
rect 14096 10406 14148 10412
rect 14108 10062 14136 10406
rect 14096 10056 14148 10062
rect 14096 9998 14148 10004
rect 13820 8628 13872 8634
rect 13820 8570 13872 8576
rect 14004 8628 14056 8634
rect 14004 8570 14056 8576
rect 13728 8492 13780 8498
rect 13728 8434 13780 8440
rect 14096 8492 14148 8498
rect 14096 8434 14148 8440
rect 13740 6934 13768 8434
rect 14108 7954 14136 8434
rect 14096 7948 14148 7954
rect 14096 7890 14148 7896
rect 14108 7546 14136 7890
rect 14096 7540 14148 7546
rect 14096 7482 14148 7488
rect 13728 6928 13780 6934
rect 13728 6870 13780 6876
rect 13268 6792 13320 6798
rect 13268 6734 13320 6740
rect 13544 6792 13596 6798
rect 13544 6734 13596 6740
rect 12808 6724 12860 6730
rect 12808 6666 12860 6672
rect 12532 6452 12584 6458
rect 12452 6412 12532 6440
rect 12256 6394 12308 6400
rect 12532 6394 12584 6400
rect 12164 6316 12216 6322
rect 12164 6258 12216 6264
rect 12820 6118 12848 6666
rect 13280 6390 13308 6734
rect 13912 6724 13964 6730
rect 13912 6666 13964 6672
rect 14004 6724 14056 6730
rect 14004 6666 14056 6672
rect 13268 6384 13320 6390
rect 13268 6326 13320 6332
rect 11704 6112 11756 6118
rect 11704 6054 11756 6060
rect 12072 6112 12124 6118
rect 12072 6054 12124 6060
rect 12808 6112 12860 6118
rect 12808 6054 12860 6060
rect 11612 5908 11664 5914
rect 11612 5850 11664 5856
rect 11716 5642 11744 6054
rect 12820 5914 12848 6054
rect 12808 5908 12860 5914
rect 12808 5850 12860 5856
rect 13924 5778 13952 6666
rect 14016 6458 14044 6666
rect 14004 6452 14056 6458
rect 14004 6394 14056 6400
rect 14292 5778 14320 13790
rect 14556 13738 14608 13744
rect 14568 13394 14596 13738
rect 14660 13394 14688 15030
rect 14740 14408 14792 14414
rect 14740 14350 14792 14356
rect 14752 14074 14780 14350
rect 14740 14068 14792 14074
rect 14740 14010 14792 14016
rect 14844 13530 14872 16680
rect 14936 13802 14964 17682
rect 15028 17542 15056 18294
rect 15016 17536 15068 17542
rect 15016 17478 15068 17484
rect 15212 17270 15240 22374
rect 15304 21146 15332 22918
rect 15580 22778 15608 22986
rect 15568 22772 15620 22778
rect 15568 22714 15620 22720
rect 15568 22636 15620 22642
rect 15568 22578 15620 22584
rect 15580 22166 15608 22578
rect 15568 22160 15620 22166
rect 15568 22102 15620 22108
rect 15292 21140 15344 21146
rect 15292 21082 15344 21088
rect 15292 19168 15344 19174
rect 15292 19110 15344 19116
rect 15304 17814 15332 19110
rect 15384 18964 15436 18970
rect 15384 18906 15436 18912
rect 15396 17882 15424 18906
rect 15672 18222 15700 24346
rect 16304 24268 16356 24274
rect 16304 24210 16356 24216
rect 16316 23866 16344 24210
rect 16920 23964 17296 23973
rect 16976 23962 17000 23964
rect 17056 23962 17080 23964
rect 17136 23962 17160 23964
rect 17216 23962 17240 23964
rect 16976 23910 16986 23962
rect 17230 23910 17240 23962
rect 16976 23908 17000 23910
rect 17056 23908 17080 23910
rect 17136 23908 17160 23910
rect 17216 23908 17240 23910
rect 16920 23899 17296 23908
rect 16028 23860 16080 23866
rect 16028 23802 16080 23808
rect 16304 23860 16356 23866
rect 16304 23802 16356 23808
rect 15936 23248 15988 23254
rect 15936 23190 15988 23196
rect 15752 23112 15804 23118
rect 15752 23054 15804 23060
rect 15764 22098 15792 23054
rect 15844 22976 15896 22982
rect 15844 22918 15896 22924
rect 15856 22778 15884 22918
rect 15844 22772 15896 22778
rect 15844 22714 15896 22720
rect 15948 22574 15976 23190
rect 16040 22642 16068 23802
rect 16180 23420 16556 23429
rect 16236 23418 16260 23420
rect 16316 23418 16340 23420
rect 16396 23418 16420 23420
rect 16476 23418 16500 23420
rect 16236 23366 16246 23418
rect 16490 23366 16500 23418
rect 16236 23364 16260 23366
rect 16316 23364 16340 23366
rect 16396 23364 16420 23366
rect 16476 23364 16500 23366
rect 16180 23355 16556 23364
rect 16212 23044 16264 23050
rect 16212 22986 16264 22992
rect 17592 23044 17644 23050
rect 17592 22986 17644 22992
rect 16224 22778 16252 22986
rect 16920 22876 17296 22885
rect 16976 22874 17000 22876
rect 17056 22874 17080 22876
rect 17136 22874 17160 22876
rect 17216 22874 17240 22876
rect 16976 22822 16986 22874
rect 17230 22822 17240 22874
rect 16976 22820 17000 22822
rect 17056 22820 17080 22822
rect 17136 22820 17160 22822
rect 17216 22820 17240 22822
rect 16920 22811 17296 22820
rect 16212 22772 16264 22778
rect 16212 22714 16264 22720
rect 16028 22636 16080 22642
rect 16028 22578 16080 22584
rect 15936 22568 15988 22574
rect 15936 22510 15988 22516
rect 15844 22432 15896 22438
rect 15844 22374 15896 22380
rect 15856 22098 15884 22374
rect 15752 22092 15804 22098
rect 15752 22034 15804 22040
rect 15844 22092 15896 22098
rect 15948 22094 15976 22510
rect 16180 22332 16556 22341
rect 16236 22330 16260 22332
rect 16316 22330 16340 22332
rect 16396 22330 16420 22332
rect 16476 22330 16500 22332
rect 16236 22278 16246 22330
rect 16490 22278 16500 22330
rect 16236 22276 16260 22278
rect 16316 22276 16340 22278
rect 16396 22276 16420 22278
rect 16476 22276 16500 22278
rect 16180 22267 16556 22276
rect 15948 22066 16160 22094
rect 15844 22034 15896 22040
rect 16132 22030 16160 22066
rect 16120 22024 16172 22030
rect 16120 21966 16172 21972
rect 17316 21888 17368 21894
rect 17316 21830 17368 21836
rect 16920 21788 17296 21797
rect 16976 21786 17000 21788
rect 17056 21786 17080 21788
rect 17136 21786 17160 21788
rect 17216 21786 17240 21788
rect 16976 21734 16986 21786
rect 17230 21734 17240 21786
rect 16976 21732 17000 21734
rect 17056 21732 17080 21734
rect 17136 21732 17160 21734
rect 17216 21732 17240 21734
rect 16920 21723 17296 21732
rect 17328 21350 17356 21830
rect 17604 21690 17632 22986
rect 17972 22778 18000 24686
rect 18236 23588 18288 23594
rect 18236 23530 18288 23536
rect 18248 23118 18276 23530
rect 18236 23112 18288 23118
rect 18236 23054 18288 23060
rect 17960 22772 18012 22778
rect 17960 22714 18012 22720
rect 18340 22094 18368 26250
rect 18524 25294 18552 27406
rect 18604 27328 18656 27334
rect 18604 27270 18656 27276
rect 18696 27328 18748 27334
rect 18696 27270 18748 27276
rect 18616 26586 18644 27270
rect 18708 27130 18736 27270
rect 18696 27124 18748 27130
rect 18696 27066 18748 27072
rect 18696 26784 18748 26790
rect 18696 26726 18748 26732
rect 18788 26784 18840 26790
rect 18788 26726 18840 26732
rect 18708 26586 18736 26726
rect 18604 26580 18656 26586
rect 18604 26522 18656 26528
rect 18696 26580 18748 26586
rect 18696 26522 18748 26528
rect 18800 26246 18828 26726
rect 18788 26240 18840 26246
rect 18788 26182 18840 26188
rect 18512 25288 18564 25294
rect 18512 25230 18564 25236
rect 18420 24744 18472 24750
rect 18420 24686 18472 24692
rect 18432 24410 18460 24686
rect 18892 24410 18920 28018
rect 18972 28008 19024 28014
rect 18972 27950 19024 27956
rect 18984 27470 19012 27950
rect 19352 27538 19380 30670
rect 19444 29850 19472 31350
rect 20180 31210 20208 31758
rect 22920 31580 23296 31589
rect 22976 31578 23000 31580
rect 23056 31578 23080 31580
rect 23136 31578 23160 31580
rect 23216 31578 23240 31580
rect 22976 31526 22986 31578
rect 23230 31526 23240 31578
rect 22976 31524 23000 31526
rect 23056 31524 23080 31526
rect 23136 31524 23160 31526
rect 23216 31524 23240 31526
rect 22920 31515 23296 31524
rect 24688 31482 24716 32370
rect 30564 32224 30616 32230
rect 30564 32166 30616 32172
rect 28180 32124 28556 32133
rect 28236 32122 28260 32124
rect 28316 32122 28340 32124
rect 28396 32122 28420 32124
rect 28476 32122 28500 32124
rect 28236 32070 28246 32122
rect 28490 32070 28500 32122
rect 28236 32068 28260 32070
rect 28316 32068 28340 32070
rect 28396 32068 28420 32070
rect 28476 32068 28500 32070
rect 28180 32059 28556 32068
rect 28920 31580 29296 31589
rect 28976 31578 29000 31580
rect 29056 31578 29080 31580
rect 29136 31578 29160 31580
rect 29216 31578 29240 31580
rect 28976 31526 28986 31578
rect 29230 31526 29240 31578
rect 28976 31524 29000 31526
rect 29056 31524 29080 31526
rect 29136 31524 29160 31526
rect 29216 31524 29240 31526
rect 28920 31515 29296 31524
rect 24676 31476 24728 31482
rect 24676 31418 24728 31424
rect 20168 31204 20220 31210
rect 20168 31146 20220 31152
rect 19524 30660 19576 30666
rect 19524 30602 19576 30608
rect 19536 30190 19564 30602
rect 19708 30320 19760 30326
rect 19708 30262 19760 30268
rect 19524 30184 19576 30190
rect 19524 30126 19576 30132
rect 19720 29850 19748 30262
rect 19432 29844 19484 29850
rect 19432 29786 19484 29792
rect 19708 29844 19760 29850
rect 19708 29786 19760 29792
rect 20180 28014 20208 31146
rect 22180 31036 22556 31045
rect 22236 31034 22260 31036
rect 22316 31034 22340 31036
rect 22396 31034 22420 31036
rect 22476 31034 22500 31036
rect 22236 30982 22246 31034
rect 22490 30982 22500 31034
rect 22236 30980 22260 30982
rect 22316 30980 22340 30982
rect 22396 30980 22420 30982
rect 22476 30980 22500 30982
rect 22180 30971 22556 30980
rect 28180 31036 28556 31045
rect 28236 31034 28260 31036
rect 28316 31034 28340 31036
rect 28396 31034 28420 31036
rect 28476 31034 28500 31036
rect 28236 30982 28246 31034
rect 28490 30982 28500 31034
rect 28236 30980 28260 30982
rect 28316 30980 28340 30982
rect 28396 30980 28420 30982
rect 28476 30980 28500 30982
rect 28180 30971 28556 30980
rect 22920 30492 23296 30501
rect 22976 30490 23000 30492
rect 23056 30490 23080 30492
rect 23136 30490 23160 30492
rect 23216 30490 23240 30492
rect 22976 30438 22986 30490
rect 23230 30438 23240 30490
rect 22976 30436 23000 30438
rect 23056 30436 23080 30438
rect 23136 30436 23160 30438
rect 23216 30436 23240 30438
rect 22920 30427 23296 30436
rect 28920 30492 29296 30501
rect 28976 30490 29000 30492
rect 29056 30490 29080 30492
rect 29136 30490 29160 30492
rect 29216 30490 29240 30492
rect 28976 30438 28986 30490
rect 29230 30438 29240 30490
rect 28976 30436 29000 30438
rect 29056 30436 29080 30438
rect 29136 30436 29160 30438
rect 29216 30436 29240 30438
rect 28920 30427 29296 30436
rect 20444 30048 20496 30054
rect 20444 29990 20496 29996
rect 20456 29646 20484 29990
rect 22180 29948 22556 29957
rect 22236 29946 22260 29948
rect 22316 29946 22340 29948
rect 22396 29946 22420 29948
rect 22476 29946 22500 29948
rect 22236 29894 22246 29946
rect 22490 29894 22500 29946
rect 22236 29892 22260 29894
rect 22316 29892 22340 29894
rect 22396 29892 22420 29894
rect 22476 29892 22500 29894
rect 22180 29883 22556 29892
rect 28180 29948 28556 29957
rect 28236 29946 28260 29948
rect 28316 29946 28340 29948
rect 28396 29946 28420 29948
rect 28476 29946 28500 29948
rect 28236 29894 28246 29946
rect 28490 29894 28500 29946
rect 28236 29892 28260 29894
rect 28316 29892 28340 29894
rect 28396 29892 28420 29894
rect 28476 29892 28500 29894
rect 28180 29883 28556 29892
rect 20444 29640 20496 29646
rect 20444 29582 20496 29588
rect 20352 28076 20404 28082
rect 20352 28018 20404 28024
rect 20168 28008 20220 28014
rect 20168 27950 20220 27956
rect 19984 27940 20036 27946
rect 19984 27882 20036 27888
rect 19708 27600 19760 27606
rect 19708 27542 19760 27548
rect 19340 27532 19392 27538
rect 19340 27474 19392 27480
rect 18972 27464 19024 27470
rect 18972 27406 19024 27412
rect 19156 26920 19208 26926
rect 19156 26862 19208 26868
rect 19168 26586 19196 26862
rect 19340 26852 19392 26858
rect 19340 26794 19392 26800
rect 19156 26580 19208 26586
rect 19156 26522 19208 26528
rect 18420 24404 18472 24410
rect 18420 24346 18472 24352
rect 18880 24404 18932 24410
rect 18880 24346 18932 24352
rect 19064 24200 19116 24206
rect 19064 24142 19116 24148
rect 18880 23588 18932 23594
rect 18880 23530 18932 23536
rect 18420 23316 18472 23322
rect 18420 23258 18472 23264
rect 18432 23050 18460 23258
rect 18892 23118 18920 23530
rect 18604 23112 18656 23118
rect 18604 23054 18656 23060
rect 18880 23112 18932 23118
rect 18880 23054 18932 23060
rect 18420 23044 18472 23050
rect 18420 22986 18472 22992
rect 18512 22976 18564 22982
rect 18512 22918 18564 22924
rect 18248 22066 18368 22094
rect 17592 21684 17644 21690
rect 17592 21626 17644 21632
rect 17316 21344 17368 21350
rect 17316 21286 17368 21292
rect 16180 21244 16556 21253
rect 16236 21242 16260 21244
rect 16316 21242 16340 21244
rect 16396 21242 16420 21244
rect 16476 21242 16500 21244
rect 16236 21190 16246 21242
rect 16490 21190 16500 21242
rect 16236 21188 16260 21190
rect 16316 21188 16340 21190
rect 16396 21188 16420 21190
rect 16476 21188 16500 21190
rect 16180 21179 16556 21188
rect 16920 20700 17296 20709
rect 16976 20698 17000 20700
rect 17056 20698 17080 20700
rect 17136 20698 17160 20700
rect 17216 20698 17240 20700
rect 16976 20646 16986 20698
rect 17230 20646 17240 20698
rect 16976 20644 17000 20646
rect 17056 20644 17080 20646
rect 17136 20644 17160 20646
rect 17216 20644 17240 20646
rect 16920 20635 17296 20644
rect 16180 20156 16556 20165
rect 16236 20154 16260 20156
rect 16316 20154 16340 20156
rect 16396 20154 16420 20156
rect 16476 20154 16500 20156
rect 16236 20102 16246 20154
rect 16490 20102 16500 20154
rect 16236 20100 16260 20102
rect 16316 20100 16340 20102
rect 16396 20100 16420 20102
rect 16476 20100 16500 20102
rect 16180 20091 16556 20100
rect 17684 19848 17736 19854
rect 17684 19790 17736 19796
rect 17500 19712 17552 19718
rect 17500 19654 17552 19660
rect 16920 19612 17296 19621
rect 16976 19610 17000 19612
rect 17056 19610 17080 19612
rect 17136 19610 17160 19612
rect 17216 19610 17240 19612
rect 16976 19558 16986 19610
rect 17230 19558 17240 19610
rect 16976 19556 17000 19558
rect 17056 19556 17080 19558
rect 17136 19556 17160 19558
rect 17216 19556 17240 19558
rect 16920 19547 17296 19556
rect 17512 19446 17540 19654
rect 15936 19440 15988 19446
rect 15936 19382 15988 19388
rect 17500 19440 17552 19446
rect 17500 19382 17552 19388
rect 15948 18970 15976 19382
rect 17316 19372 17368 19378
rect 17316 19314 17368 19320
rect 16180 19068 16556 19077
rect 16236 19066 16260 19068
rect 16316 19066 16340 19068
rect 16396 19066 16420 19068
rect 16476 19066 16500 19068
rect 16236 19014 16246 19066
rect 16490 19014 16500 19066
rect 16236 19012 16260 19014
rect 16316 19012 16340 19014
rect 16396 19012 16420 19014
rect 16476 19012 16500 19014
rect 16180 19003 16556 19012
rect 15936 18964 15988 18970
rect 15936 18906 15988 18912
rect 16672 18896 16724 18902
rect 16672 18838 16724 18844
rect 16212 18624 16264 18630
rect 16212 18566 16264 18572
rect 16224 18426 16252 18566
rect 16684 18426 16712 18838
rect 16920 18524 17296 18533
rect 16976 18522 17000 18524
rect 17056 18522 17080 18524
rect 17136 18522 17160 18524
rect 17216 18522 17240 18524
rect 16976 18470 16986 18522
rect 17230 18470 17240 18522
rect 16976 18468 17000 18470
rect 17056 18468 17080 18470
rect 17136 18468 17160 18470
rect 17216 18468 17240 18470
rect 16920 18459 17296 18468
rect 16212 18420 16264 18426
rect 16212 18362 16264 18368
rect 16672 18420 16724 18426
rect 16672 18362 16724 18368
rect 17328 18290 17356 19314
rect 17696 18970 17724 19790
rect 17684 18964 17736 18970
rect 17684 18906 17736 18912
rect 18248 18834 18276 22066
rect 18524 22030 18552 22918
rect 18616 22506 18644 23054
rect 19076 22642 19104 24142
rect 19064 22636 19116 22642
rect 19064 22578 19116 22584
rect 18604 22500 18656 22506
rect 18604 22442 18656 22448
rect 18512 22024 18564 22030
rect 18512 21966 18564 21972
rect 18616 21554 18644 22442
rect 19076 22094 19104 22578
rect 18892 22066 19104 22094
rect 18604 21548 18656 21554
rect 18604 21490 18656 21496
rect 18328 19712 18380 19718
rect 18328 19654 18380 19660
rect 18236 18828 18288 18834
rect 17972 18788 18236 18816
rect 17316 18284 17368 18290
rect 17316 18226 17368 18232
rect 15660 18216 15712 18222
rect 15660 18158 15712 18164
rect 15384 17876 15436 17882
rect 15384 17818 15436 17824
rect 15292 17808 15344 17814
rect 15292 17750 15344 17756
rect 15476 17740 15528 17746
rect 15476 17682 15528 17688
rect 15200 17264 15252 17270
rect 15200 17206 15252 17212
rect 15200 16788 15252 16794
rect 15200 16730 15252 16736
rect 15212 16114 15240 16730
rect 15200 16108 15252 16114
rect 15200 16050 15252 16056
rect 15384 13864 15436 13870
rect 15384 13806 15436 13812
rect 14924 13796 14976 13802
rect 14924 13738 14976 13744
rect 14832 13524 14884 13530
rect 14832 13466 14884 13472
rect 14556 13388 14608 13394
rect 14556 13330 14608 13336
rect 14648 13388 14700 13394
rect 14700 13348 14780 13376
rect 14648 13330 14700 13336
rect 14372 12844 14424 12850
rect 14372 12786 14424 12792
rect 14384 8838 14412 12786
rect 14648 9920 14700 9926
rect 14648 9862 14700 9868
rect 14660 9654 14688 9862
rect 14648 9648 14700 9654
rect 14648 9590 14700 9596
rect 14372 8832 14424 8838
rect 14372 8774 14424 8780
rect 14384 8498 14412 8774
rect 14372 8492 14424 8498
rect 14372 8434 14424 8440
rect 14556 8492 14608 8498
rect 14556 8434 14608 8440
rect 13912 5772 13964 5778
rect 13912 5714 13964 5720
rect 14280 5772 14332 5778
rect 14280 5714 14332 5720
rect 12164 5704 12216 5710
rect 12164 5646 12216 5652
rect 12808 5704 12860 5710
rect 12808 5646 12860 5652
rect 11704 5636 11756 5642
rect 11704 5578 11756 5584
rect 10920 5468 11296 5477
rect 10976 5466 11000 5468
rect 11056 5466 11080 5468
rect 11136 5466 11160 5468
rect 11216 5466 11240 5468
rect 10976 5414 10986 5466
rect 11230 5414 11240 5466
rect 10976 5412 11000 5414
rect 11056 5412 11080 5414
rect 11136 5412 11160 5414
rect 11216 5412 11240 5414
rect 10920 5403 11296 5412
rect 10704 4678 10824 4706
rect 10600 4140 10652 4146
rect 10600 4082 10652 4088
rect 10704 4078 10732 4678
rect 10784 4616 10836 4622
rect 10784 4558 10836 4564
rect 10048 4072 10100 4078
rect 9692 3998 9812 4026
rect 10048 4014 10100 4020
rect 10692 4072 10744 4078
rect 10692 4014 10744 4020
rect 9680 3936 9732 3942
rect 9680 3878 9732 3884
rect 9692 3738 9720 3878
rect 9680 3732 9732 3738
rect 9680 3674 9732 3680
rect 9784 3534 9812 3998
rect 10048 3936 10100 3942
rect 10048 3878 10100 3884
rect 10060 3738 10088 3878
rect 10180 3836 10556 3845
rect 10236 3834 10260 3836
rect 10316 3834 10340 3836
rect 10396 3834 10420 3836
rect 10476 3834 10500 3836
rect 10236 3782 10246 3834
rect 10490 3782 10500 3834
rect 10236 3780 10260 3782
rect 10316 3780 10340 3782
rect 10396 3780 10420 3782
rect 10476 3780 10500 3782
rect 10180 3771 10556 3780
rect 10048 3732 10100 3738
rect 10048 3674 10100 3680
rect 9772 3528 9824 3534
rect 9772 3470 9824 3476
rect 9036 3460 9088 3466
rect 9036 3402 9088 3408
rect 9048 3058 9076 3402
rect 9496 3392 9548 3398
rect 9496 3334 9548 3340
rect 9508 3194 9536 3334
rect 9496 3188 9548 3194
rect 9496 3130 9548 3136
rect 6920 3052 6972 3058
rect 6920 2994 6972 3000
rect 9036 3052 9088 3058
rect 9036 2994 9088 3000
rect 9784 2990 9812 3470
rect 9864 3392 9916 3398
rect 9864 3334 9916 3340
rect 9876 3126 9904 3334
rect 10796 3194 10824 4558
rect 10920 4380 11296 4389
rect 10976 4378 11000 4380
rect 11056 4378 11080 4380
rect 11136 4378 11160 4380
rect 11216 4378 11240 4380
rect 10976 4326 10986 4378
rect 11230 4326 11240 4378
rect 10976 4324 11000 4326
rect 11056 4324 11080 4326
rect 11136 4324 11160 4326
rect 11216 4324 11240 4326
rect 10920 4315 11296 4324
rect 11888 4072 11940 4078
rect 11888 4014 11940 4020
rect 11612 3460 11664 3466
rect 11612 3402 11664 3408
rect 10920 3292 11296 3301
rect 10976 3290 11000 3292
rect 11056 3290 11080 3292
rect 11136 3290 11160 3292
rect 11216 3290 11240 3292
rect 10976 3238 10986 3290
rect 11230 3238 11240 3290
rect 10976 3236 11000 3238
rect 11056 3236 11080 3238
rect 11136 3236 11160 3238
rect 11216 3236 11240 3238
rect 10920 3227 11296 3236
rect 11624 3194 11652 3402
rect 11900 3398 11928 4014
rect 12176 3602 12204 5646
rect 12820 5166 12848 5646
rect 13924 5370 13952 5714
rect 14096 5568 14148 5574
rect 14096 5510 14148 5516
rect 13912 5364 13964 5370
rect 13912 5306 13964 5312
rect 13084 5228 13136 5234
rect 13084 5170 13136 5176
rect 12808 5160 12860 5166
rect 12808 5102 12860 5108
rect 13096 4826 13124 5170
rect 14108 4826 14136 5510
rect 14292 5302 14320 5714
rect 14280 5296 14332 5302
rect 14280 5238 14332 5244
rect 13084 4820 13136 4826
rect 13084 4762 13136 4768
rect 14096 4820 14148 4826
rect 14096 4762 14148 4768
rect 14568 3602 14596 8434
rect 14752 7342 14780 13348
rect 14844 10470 14872 13466
rect 14936 12434 14964 13738
rect 15396 13734 15424 13806
rect 15384 13728 15436 13734
rect 15384 13670 15436 13676
rect 15488 12434 15516 17682
rect 15568 15904 15620 15910
rect 15568 15846 15620 15852
rect 15580 15706 15608 15846
rect 15568 15700 15620 15706
rect 15568 15642 15620 15648
rect 15672 15586 15700 18158
rect 16180 17980 16556 17989
rect 16236 17978 16260 17980
rect 16316 17978 16340 17980
rect 16396 17978 16420 17980
rect 16476 17978 16500 17980
rect 16236 17926 16246 17978
rect 16490 17926 16500 17978
rect 16236 17924 16260 17926
rect 16316 17924 16340 17926
rect 16396 17924 16420 17926
rect 16476 17924 16500 17926
rect 16180 17915 16556 17924
rect 16488 17672 16540 17678
rect 16488 17614 16540 17620
rect 15844 17536 15896 17542
rect 15844 17478 15896 17484
rect 15856 17338 15884 17478
rect 16500 17338 16528 17614
rect 16920 17436 17296 17445
rect 16976 17434 17000 17436
rect 17056 17434 17080 17436
rect 17136 17434 17160 17436
rect 17216 17434 17240 17436
rect 16976 17382 16986 17434
rect 17230 17382 17240 17434
rect 16976 17380 17000 17382
rect 17056 17380 17080 17382
rect 17136 17380 17160 17382
rect 17216 17380 17240 17382
rect 16920 17371 17296 17380
rect 15844 17332 15896 17338
rect 15844 17274 15896 17280
rect 16488 17332 16540 17338
rect 16488 17274 16540 17280
rect 15752 17264 15804 17270
rect 15752 17206 15804 17212
rect 15764 16114 15792 17206
rect 17328 17202 17356 18226
rect 17868 17536 17920 17542
rect 17866 17504 17868 17513
rect 17920 17504 17922 17513
rect 17866 17439 17922 17448
rect 17316 17196 17368 17202
rect 17316 17138 17368 17144
rect 16180 16892 16556 16901
rect 16236 16890 16260 16892
rect 16316 16890 16340 16892
rect 16396 16890 16420 16892
rect 16476 16890 16500 16892
rect 16236 16838 16246 16890
rect 16490 16838 16500 16890
rect 16236 16836 16260 16838
rect 16316 16836 16340 16838
rect 16396 16836 16420 16838
rect 16476 16836 16500 16838
rect 16180 16827 16556 16836
rect 16920 16348 17296 16357
rect 16976 16346 17000 16348
rect 17056 16346 17080 16348
rect 17136 16346 17160 16348
rect 17216 16346 17240 16348
rect 16976 16294 16986 16346
rect 17230 16294 17240 16346
rect 16976 16292 17000 16294
rect 17056 16292 17080 16294
rect 17136 16292 17160 16294
rect 17216 16292 17240 16294
rect 16920 16283 17296 16292
rect 15752 16108 15804 16114
rect 15752 16050 15804 16056
rect 14936 12406 15056 12434
rect 14832 10464 14884 10470
rect 14832 10406 14884 10412
rect 14832 10056 14884 10062
rect 14832 9998 14884 10004
rect 14844 9178 14872 9998
rect 14924 9988 14976 9994
rect 14924 9930 14976 9936
rect 14832 9172 14884 9178
rect 14832 9114 14884 9120
rect 14830 8528 14886 8537
rect 14936 8498 14964 9930
rect 15028 9042 15056 12406
rect 15396 12406 15516 12434
rect 15580 15558 15700 15586
rect 15292 12300 15344 12306
rect 15292 12242 15344 12248
rect 15108 10668 15160 10674
rect 15108 10610 15160 10616
rect 15016 9036 15068 9042
rect 15016 8978 15068 8984
rect 15120 8838 15148 10610
rect 15304 10606 15332 12242
rect 15292 10600 15344 10606
rect 15292 10542 15344 10548
rect 15396 9466 15424 12406
rect 15580 12306 15608 15558
rect 15764 13938 15792 16050
rect 17972 15910 18000 18788
rect 18236 18770 18288 18776
rect 18340 18766 18368 19654
rect 18328 18760 18380 18766
rect 18328 18702 18380 18708
rect 18052 18692 18104 18698
rect 18052 18634 18104 18640
rect 18064 18426 18092 18634
rect 18052 18420 18104 18426
rect 18052 18362 18104 18368
rect 18418 17640 18474 17649
rect 18418 17575 18420 17584
rect 18472 17575 18474 17584
rect 18420 17546 18472 17552
rect 18236 17196 18288 17202
rect 18236 17138 18288 17144
rect 18248 16794 18276 17138
rect 18236 16788 18288 16794
rect 18236 16730 18288 16736
rect 17960 15904 18012 15910
rect 17960 15846 18012 15852
rect 16180 15804 16556 15813
rect 16236 15802 16260 15804
rect 16316 15802 16340 15804
rect 16396 15802 16420 15804
rect 16476 15802 16500 15804
rect 16236 15750 16246 15802
rect 16490 15750 16500 15802
rect 16236 15748 16260 15750
rect 16316 15748 16340 15750
rect 16396 15748 16420 15750
rect 16476 15748 16500 15750
rect 16180 15739 16556 15748
rect 17776 15496 17828 15502
rect 17776 15438 17828 15444
rect 17592 15360 17644 15366
rect 17592 15302 17644 15308
rect 16920 15260 17296 15269
rect 16976 15258 17000 15260
rect 17056 15258 17080 15260
rect 17136 15258 17160 15260
rect 17216 15258 17240 15260
rect 16976 15206 16986 15258
rect 17230 15206 17240 15258
rect 16976 15204 17000 15206
rect 17056 15204 17080 15206
rect 17136 15204 17160 15206
rect 17216 15204 17240 15206
rect 16920 15195 17296 15204
rect 17604 15026 17632 15302
rect 17592 15020 17644 15026
rect 17592 14962 17644 14968
rect 16180 14716 16556 14725
rect 16236 14714 16260 14716
rect 16316 14714 16340 14716
rect 16396 14714 16420 14716
rect 16476 14714 16500 14716
rect 16236 14662 16246 14714
rect 16490 14662 16500 14714
rect 16236 14660 16260 14662
rect 16316 14660 16340 14662
rect 16396 14660 16420 14662
rect 16476 14660 16500 14662
rect 16180 14651 16556 14660
rect 17788 14618 17816 15438
rect 17972 14618 18000 15846
rect 18144 15496 18196 15502
rect 18144 15438 18196 15444
rect 18236 15496 18288 15502
rect 18236 15438 18288 15444
rect 18052 15428 18104 15434
rect 18052 15370 18104 15376
rect 17776 14612 17828 14618
rect 17776 14554 17828 14560
rect 17960 14612 18012 14618
rect 17960 14554 18012 14560
rect 16028 14544 16080 14550
rect 17972 14498 18000 14554
rect 16028 14486 16080 14492
rect 16040 14006 16068 14486
rect 17880 14470 18000 14498
rect 16120 14272 16172 14278
rect 16120 14214 16172 14220
rect 16672 14272 16724 14278
rect 16672 14214 16724 14220
rect 16132 14074 16160 14214
rect 16120 14068 16172 14074
rect 16120 14010 16172 14016
rect 16028 14000 16080 14006
rect 16028 13942 16080 13948
rect 16684 13938 16712 14214
rect 16920 14172 17296 14181
rect 16976 14170 17000 14172
rect 17056 14170 17080 14172
rect 17136 14170 17160 14172
rect 17216 14170 17240 14172
rect 16976 14118 16986 14170
rect 17230 14118 17240 14170
rect 16976 14116 17000 14118
rect 17056 14116 17080 14118
rect 17136 14116 17160 14118
rect 17216 14116 17240 14118
rect 16920 14107 17296 14116
rect 15752 13932 15804 13938
rect 15752 13874 15804 13880
rect 16672 13932 16724 13938
rect 16672 13874 16724 13880
rect 15660 13184 15712 13190
rect 15660 13126 15712 13132
rect 15568 12300 15620 12306
rect 15568 12242 15620 12248
rect 15476 11008 15528 11014
rect 15476 10950 15528 10956
rect 15568 11008 15620 11014
rect 15568 10950 15620 10956
rect 15488 10130 15516 10950
rect 15580 10810 15608 10950
rect 15568 10804 15620 10810
rect 15568 10746 15620 10752
rect 15476 10124 15528 10130
rect 15476 10066 15528 10072
rect 15304 9438 15424 9466
rect 15108 8832 15160 8838
rect 15108 8774 15160 8780
rect 14830 8463 14832 8472
rect 14884 8463 14886 8472
rect 14924 8492 14976 8498
rect 14832 8434 14884 8440
rect 14924 8434 14976 8440
rect 15120 7342 15148 8774
rect 14740 7336 14792 7342
rect 14740 7278 14792 7284
rect 15108 7336 15160 7342
rect 15108 7278 15160 7284
rect 14648 7200 14700 7206
rect 14648 7142 14700 7148
rect 14660 6458 14688 7142
rect 14648 6452 14700 6458
rect 14648 6394 14700 6400
rect 15120 5574 15148 7278
rect 15108 5568 15160 5574
rect 15108 5510 15160 5516
rect 15200 4684 15252 4690
rect 15200 4626 15252 4632
rect 15016 4480 15068 4486
rect 15016 4422 15068 4428
rect 15028 4282 15056 4422
rect 15016 4276 15068 4282
rect 15016 4218 15068 4224
rect 14648 4004 14700 4010
rect 14648 3946 14700 3952
rect 14660 3602 14688 3946
rect 15212 3670 15240 4626
rect 15304 4146 15332 9438
rect 15384 9376 15436 9382
rect 15384 9318 15436 9324
rect 15396 9178 15424 9318
rect 15384 9172 15436 9178
rect 15384 9114 15436 9120
rect 15476 8560 15528 8566
rect 15476 8502 15528 8508
rect 15382 7304 15438 7313
rect 15488 7274 15516 8502
rect 15382 7239 15438 7248
rect 15476 7268 15528 7274
rect 15396 7002 15424 7239
rect 15476 7210 15528 7216
rect 15488 7002 15516 7210
rect 15384 6996 15436 7002
rect 15384 6938 15436 6944
rect 15476 6996 15528 7002
rect 15476 6938 15528 6944
rect 15476 5024 15528 5030
rect 15476 4966 15528 4972
rect 15488 4554 15516 4966
rect 15476 4548 15528 4554
rect 15476 4490 15528 4496
rect 15292 4140 15344 4146
rect 15292 4082 15344 4088
rect 15384 3936 15436 3942
rect 15384 3878 15436 3884
rect 15396 3738 15424 3878
rect 15384 3732 15436 3738
rect 15384 3674 15436 3680
rect 15200 3664 15252 3670
rect 15200 3606 15252 3612
rect 15488 3602 15516 4490
rect 15672 4146 15700 13126
rect 15764 9654 15792 13874
rect 16580 13864 16632 13870
rect 16580 13806 16632 13812
rect 15844 13728 15896 13734
rect 15844 13670 15896 13676
rect 16028 13728 16080 13734
rect 16028 13670 16080 13676
rect 15856 12306 15884 13670
rect 16040 13410 16068 13670
rect 16180 13628 16556 13637
rect 16236 13626 16260 13628
rect 16316 13626 16340 13628
rect 16396 13626 16420 13628
rect 16476 13626 16500 13628
rect 16236 13574 16246 13626
rect 16490 13574 16500 13626
rect 16236 13572 16260 13574
rect 16316 13572 16340 13574
rect 16396 13572 16420 13574
rect 16476 13572 16500 13574
rect 16180 13563 16556 13572
rect 16212 13524 16264 13530
rect 16212 13466 16264 13472
rect 16040 13382 16160 13410
rect 16132 13326 16160 13382
rect 16224 13326 16252 13466
rect 16592 13326 16620 13806
rect 16028 13320 16080 13326
rect 15948 13268 16028 13274
rect 15948 13262 16080 13268
rect 16120 13320 16172 13326
rect 16120 13262 16172 13268
rect 16212 13320 16264 13326
rect 16212 13262 16264 13268
rect 16580 13320 16632 13326
rect 16580 13262 16632 13268
rect 15948 13246 16068 13262
rect 15948 12986 15976 13246
rect 16028 13184 16080 13190
rect 16028 13126 16080 13132
rect 15936 12980 15988 12986
rect 15936 12922 15988 12928
rect 16040 12434 16068 13126
rect 16920 13084 17296 13093
rect 16976 13082 17000 13084
rect 17056 13082 17080 13084
rect 17136 13082 17160 13084
rect 17216 13082 17240 13084
rect 16976 13030 16986 13082
rect 17230 13030 17240 13082
rect 16976 13028 17000 13030
rect 17056 13028 17080 13030
rect 17136 13028 17160 13030
rect 17216 13028 17240 13030
rect 16920 13019 17296 13028
rect 16180 12540 16556 12549
rect 16236 12538 16260 12540
rect 16316 12538 16340 12540
rect 16396 12538 16420 12540
rect 16476 12538 16500 12540
rect 16236 12486 16246 12538
rect 16490 12486 16500 12538
rect 16236 12484 16260 12486
rect 16316 12484 16340 12486
rect 16396 12484 16420 12486
rect 16476 12484 16500 12486
rect 16180 12475 16556 12484
rect 16040 12406 16160 12434
rect 15844 12300 15896 12306
rect 15844 12242 15896 12248
rect 16132 12238 16160 12406
rect 16120 12232 16172 12238
rect 16120 12174 16172 12180
rect 16028 12096 16080 12102
rect 16028 12038 16080 12044
rect 15936 11756 15988 11762
rect 15936 11698 15988 11704
rect 15948 11234 15976 11698
rect 16040 11354 16068 12038
rect 16132 11898 16160 12174
rect 16920 11996 17296 12005
rect 16976 11994 17000 11996
rect 17056 11994 17080 11996
rect 17136 11994 17160 11996
rect 17216 11994 17240 11996
rect 16976 11942 16986 11994
rect 17230 11942 17240 11994
rect 16976 11940 17000 11942
rect 17056 11940 17080 11942
rect 17136 11940 17160 11942
rect 17216 11940 17240 11942
rect 16920 11931 17296 11940
rect 16120 11892 16172 11898
rect 16120 11834 16172 11840
rect 16180 11452 16556 11461
rect 16236 11450 16260 11452
rect 16316 11450 16340 11452
rect 16396 11450 16420 11452
rect 16476 11450 16500 11452
rect 16236 11398 16246 11450
rect 16490 11398 16500 11450
rect 16236 11396 16260 11398
rect 16316 11396 16340 11398
rect 16396 11396 16420 11398
rect 16476 11396 16500 11398
rect 16180 11387 16556 11396
rect 16028 11348 16080 11354
rect 16028 11290 16080 11296
rect 16120 11280 16172 11286
rect 15948 11228 16120 11234
rect 15948 11222 16172 11228
rect 15948 11206 16160 11222
rect 16920 10908 17296 10917
rect 16976 10906 17000 10908
rect 17056 10906 17080 10908
rect 17136 10906 17160 10908
rect 17216 10906 17240 10908
rect 16976 10854 16986 10906
rect 17230 10854 17240 10906
rect 16976 10852 17000 10854
rect 17056 10852 17080 10854
rect 17136 10852 17160 10854
rect 17216 10852 17240 10854
rect 16920 10843 17296 10852
rect 16180 10364 16556 10373
rect 16236 10362 16260 10364
rect 16316 10362 16340 10364
rect 16396 10362 16420 10364
rect 16476 10362 16500 10364
rect 16236 10310 16246 10362
rect 16490 10310 16500 10362
rect 16236 10308 16260 10310
rect 16316 10308 16340 10310
rect 16396 10308 16420 10310
rect 16476 10308 16500 10310
rect 16180 10299 16556 10308
rect 16920 9820 17296 9829
rect 16976 9818 17000 9820
rect 17056 9818 17080 9820
rect 17136 9818 17160 9820
rect 17216 9818 17240 9820
rect 16976 9766 16986 9818
rect 17230 9766 17240 9818
rect 16976 9764 17000 9766
rect 17056 9764 17080 9766
rect 17136 9764 17160 9766
rect 17216 9764 17240 9766
rect 16920 9755 17296 9764
rect 15752 9648 15804 9654
rect 15752 9590 15804 9596
rect 15752 9376 15804 9382
rect 15752 9318 15804 9324
rect 15764 8634 15792 9318
rect 16180 9276 16556 9285
rect 16236 9274 16260 9276
rect 16316 9274 16340 9276
rect 16396 9274 16420 9276
rect 16476 9274 16500 9276
rect 16236 9222 16246 9274
rect 16490 9222 16500 9274
rect 16236 9220 16260 9222
rect 16316 9220 16340 9222
rect 16396 9220 16420 9222
rect 16476 9220 16500 9222
rect 16180 9211 16556 9220
rect 16488 8832 16540 8838
rect 16488 8774 16540 8780
rect 17684 8832 17736 8838
rect 17684 8774 17736 8780
rect 16500 8634 16528 8774
rect 16920 8732 17296 8741
rect 16976 8730 17000 8732
rect 17056 8730 17080 8732
rect 17136 8730 17160 8732
rect 17216 8730 17240 8732
rect 16976 8678 16986 8730
rect 17230 8678 17240 8730
rect 16976 8676 17000 8678
rect 17056 8676 17080 8678
rect 17136 8676 17160 8678
rect 17216 8676 17240 8678
rect 16920 8667 17296 8676
rect 15752 8628 15804 8634
rect 15752 8570 15804 8576
rect 16488 8628 16540 8634
rect 16488 8570 16540 8576
rect 16672 8492 16724 8498
rect 16672 8434 16724 8440
rect 16180 8188 16556 8197
rect 16236 8186 16260 8188
rect 16316 8186 16340 8188
rect 16396 8186 16420 8188
rect 16476 8186 16500 8188
rect 16236 8134 16246 8186
rect 16490 8134 16500 8186
rect 16236 8132 16260 8134
rect 16316 8132 16340 8134
rect 16396 8132 16420 8134
rect 16476 8132 16500 8134
rect 16180 8123 16556 8132
rect 16684 7886 16712 8434
rect 16856 8288 16908 8294
rect 16856 8230 16908 8236
rect 17316 8288 17368 8294
rect 17316 8230 17368 8236
rect 16868 7886 16896 8230
rect 16672 7880 16724 7886
rect 16672 7822 16724 7828
rect 16856 7880 16908 7886
rect 16856 7822 16908 7828
rect 16580 7744 16632 7750
rect 16580 7686 16632 7692
rect 16180 7100 16556 7109
rect 16236 7098 16260 7100
rect 16316 7098 16340 7100
rect 16396 7098 16420 7100
rect 16476 7098 16500 7100
rect 16236 7046 16246 7098
rect 16490 7046 16500 7098
rect 16236 7044 16260 7046
rect 16316 7044 16340 7046
rect 16396 7044 16420 7046
rect 16476 7044 16500 7046
rect 16180 7035 16556 7044
rect 16592 7002 16620 7686
rect 16580 6996 16632 7002
rect 16580 6938 16632 6944
rect 16684 6866 16712 7822
rect 16920 7644 17296 7653
rect 16976 7642 17000 7644
rect 17056 7642 17080 7644
rect 17136 7642 17160 7644
rect 17216 7642 17240 7644
rect 16976 7590 16986 7642
rect 17230 7590 17240 7642
rect 16976 7588 17000 7590
rect 17056 7588 17080 7590
rect 17136 7588 17160 7590
rect 17216 7588 17240 7590
rect 16920 7579 17296 7588
rect 16672 6860 16724 6866
rect 16672 6802 16724 6808
rect 16180 6012 16556 6021
rect 16236 6010 16260 6012
rect 16316 6010 16340 6012
rect 16396 6010 16420 6012
rect 16476 6010 16500 6012
rect 16236 5958 16246 6010
rect 16490 5958 16500 6010
rect 16236 5956 16260 5958
rect 16316 5956 16340 5958
rect 16396 5956 16420 5958
rect 16476 5956 16500 5958
rect 16180 5947 16556 5956
rect 16684 5778 16712 6802
rect 17328 6769 17356 8230
rect 17696 6798 17724 8774
rect 17684 6792 17736 6798
rect 17314 6760 17370 6769
rect 17684 6734 17736 6740
rect 17314 6695 17370 6704
rect 17328 6662 17356 6695
rect 16764 6656 16816 6662
rect 16764 6598 16816 6604
rect 17316 6656 17368 6662
rect 17316 6598 17368 6604
rect 16776 6254 16804 6598
rect 16920 6556 17296 6565
rect 16976 6554 17000 6556
rect 17056 6554 17080 6556
rect 17136 6554 17160 6556
rect 17216 6554 17240 6556
rect 16976 6502 16986 6554
rect 17230 6502 17240 6554
rect 16976 6500 17000 6502
rect 17056 6500 17080 6502
rect 17136 6500 17160 6502
rect 17216 6500 17240 6502
rect 16920 6491 17296 6500
rect 17696 6458 17724 6734
rect 17684 6452 17736 6458
rect 17684 6394 17736 6400
rect 17880 6254 17908 14470
rect 18064 14278 18092 15370
rect 18156 14618 18184 15438
rect 18144 14612 18196 14618
rect 18144 14554 18196 14560
rect 18248 14414 18276 15438
rect 18512 15360 18564 15366
rect 18512 15302 18564 15308
rect 18604 15360 18656 15366
rect 18604 15302 18656 15308
rect 18328 15088 18380 15094
rect 18328 15030 18380 15036
rect 18144 14408 18196 14414
rect 18144 14350 18196 14356
rect 18236 14408 18288 14414
rect 18236 14350 18288 14356
rect 18052 14272 18104 14278
rect 18052 14214 18104 14220
rect 18156 13530 18184 14350
rect 18340 14074 18368 15030
rect 18524 15026 18552 15302
rect 18512 15020 18564 15026
rect 18512 14962 18564 14968
rect 18512 14476 18564 14482
rect 18512 14418 18564 14424
rect 18328 14068 18380 14074
rect 18328 14010 18380 14016
rect 18144 13524 18196 13530
rect 18144 13466 18196 13472
rect 17960 11756 18012 11762
rect 17960 11698 18012 11704
rect 17972 11354 18000 11698
rect 17960 11348 18012 11354
rect 17960 11290 18012 11296
rect 18524 9178 18552 14418
rect 18616 14006 18644 15302
rect 18892 15144 18920 22066
rect 18972 19916 19024 19922
rect 18972 19858 19024 19864
rect 18984 19514 19012 19858
rect 18972 19508 19024 19514
rect 18972 19450 19024 19456
rect 19064 18624 19116 18630
rect 19064 18566 19116 18572
rect 19076 18426 19104 18566
rect 19064 18420 19116 18426
rect 19064 18362 19116 18368
rect 19168 18222 19196 26522
rect 19352 25974 19380 26794
rect 19720 26246 19748 27542
rect 19996 27538 20024 27882
rect 19984 27532 20036 27538
rect 19984 27474 20036 27480
rect 19892 27464 19944 27470
rect 19892 27406 19944 27412
rect 20076 27464 20128 27470
rect 20076 27406 20128 27412
rect 19708 26240 19760 26246
rect 19708 26182 19760 26188
rect 19340 25968 19392 25974
rect 19340 25910 19392 25916
rect 19904 25294 19932 27406
rect 19340 25288 19392 25294
rect 19340 25230 19392 25236
rect 19892 25288 19944 25294
rect 19892 25230 19944 25236
rect 19352 22710 19380 25230
rect 19432 25152 19484 25158
rect 19432 25094 19484 25100
rect 19444 24886 19472 25094
rect 19904 24954 19932 25230
rect 19892 24948 19944 24954
rect 20088 24936 20116 27406
rect 20260 26308 20312 26314
rect 20260 26250 20312 26256
rect 20168 26240 20220 26246
rect 20168 26182 20220 26188
rect 20180 25498 20208 26182
rect 20168 25492 20220 25498
rect 20168 25434 20220 25440
rect 19892 24890 19944 24896
rect 19996 24908 20116 24936
rect 19432 24880 19484 24886
rect 19432 24822 19484 24828
rect 19432 24608 19484 24614
rect 19432 24550 19484 24556
rect 19444 23322 19472 24550
rect 19616 24268 19668 24274
rect 19616 24210 19668 24216
rect 19524 24200 19576 24206
rect 19524 24142 19576 24148
rect 19536 23594 19564 24142
rect 19628 23798 19656 24210
rect 19996 24188 20024 24908
rect 20076 24812 20128 24818
rect 20076 24754 20128 24760
rect 20088 24410 20116 24754
rect 20076 24404 20128 24410
rect 20076 24346 20128 24352
rect 20076 24200 20128 24206
rect 19996 24160 20076 24188
rect 20076 24142 20128 24148
rect 19708 24064 19760 24070
rect 19708 24006 19760 24012
rect 19984 24064 20036 24070
rect 19984 24006 20036 24012
rect 19720 23798 19748 24006
rect 19616 23792 19668 23798
rect 19616 23734 19668 23740
rect 19708 23792 19760 23798
rect 19708 23734 19760 23740
rect 19524 23588 19576 23594
rect 19524 23530 19576 23536
rect 19432 23316 19484 23322
rect 19432 23258 19484 23264
rect 19628 23118 19656 23734
rect 19892 23724 19944 23730
rect 19892 23666 19944 23672
rect 19708 23656 19760 23662
rect 19708 23598 19760 23604
rect 19616 23112 19668 23118
rect 19616 23054 19668 23060
rect 19340 22704 19392 22710
rect 19340 22646 19392 22652
rect 19628 22642 19656 23054
rect 19616 22636 19668 22642
rect 19616 22578 19668 22584
rect 19628 22030 19656 22578
rect 19720 22094 19748 23598
rect 19904 23202 19932 23666
rect 19812 23186 19932 23202
rect 19800 23180 19932 23186
rect 19852 23174 19932 23180
rect 19800 23122 19852 23128
rect 19996 22642 20024 24006
rect 20076 23112 20128 23118
rect 20076 23054 20128 23060
rect 20088 22642 20116 23054
rect 19984 22636 20036 22642
rect 19984 22578 20036 22584
rect 20076 22636 20128 22642
rect 20076 22578 20128 22584
rect 19996 22234 20024 22578
rect 19984 22228 20036 22234
rect 19984 22170 20036 22176
rect 20180 22094 20208 25434
rect 19720 22066 19840 22094
rect 19616 22024 19668 22030
rect 19616 21966 19668 21972
rect 19340 19372 19392 19378
rect 19260 19332 19340 19360
rect 19260 18902 19288 19332
rect 19340 19314 19392 19320
rect 19708 19304 19760 19310
rect 19708 19246 19760 19252
rect 19340 19168 19392 19174
rect 19340 19110 19392 19116
rect 19248 18896 19300 18902
rect 19248 18838 19300 18844
rect 19352 18698 19380 19110
rect 19720 18986 19748 19246
rect 19628 18970 19748 18986
rect 19616 18964 19748 18970
rect 19668 18958 19748 18964
rect 19616 18906 19668 18912
rect 19340 18692 19392 18698
rect 19340 18634 19392 18640
rect 19616 18624 19668 18630
rect 19536 18572 19616 18578
rect 19536 18566 19668 18572
rect 19536 18550 19656 18566
rect 19340 18420 19392 18426
rect 19340 18362 19392 18368
rect 19156 18216 19208 18222
rect 19156 18158 19208 18164
rect 18972 18080 19024 18086
rect 18972 18022 19024 18028
rect 18984 16590 19012 18022
rect 19168 16794 19196 18158
rect 19352 17678 19380 18362
rect 19536 18154 19564 18550
rect 19720 18358 19748 18958
rect 19708 18352 19760 18358
rect 19708 18294 19760 18300
rect 19524 18148 19576 18154
rect 19524 18090 19576 18096
rect 19536 17678 19564 18090
rect 19812 17678 19840 22066
rect 20088 22066 20208 22094
rect 19984 21956 20036 21962
rect 19984 21898 20036 21904
rect 19996 19378 20024 21898
rect 19984 19372 20036 19378
rect 19984 19314 20036 19320
rect 20088 19310 20116 22066
rect 20168 19712 20220 19718
rect 20168 19654 20220 19660
rect 20180 19514 20208 19654
rect 20168 19508 20220 19514
rect 20168 19450 20220 19456
rect 20076 19304 20128 19310
rect 20076 19246 20128 19252
rect 20088 18086 20116 19246
rect 20272 18222 20300 26250
rect 20364 24290 20392 28018
rect 20456 26926 20484 29582
rect 22920 29404 23296 29413
rect 22976 29402 23000 29404
rect 23056 29402 23080 29404
rect 23136 29402 23160 29404
rect 23216 29402 23240 29404
rect 22976 29350 22986 29402
rect 23230 29350 23240 29402
rect 22976 29348 23000 29350
rect 23056 29348 23080 29350
rect 23136 29348 23160 29350
rect 23216 29348 23240 29350
rect 22920 29339 23296 29348
rect 28920 29404 29296 29413
rect 28976 29402 29000 29404
rect 29056 29402 29080 29404
rect 29136 29402 29160 29404
rect 29216 29402 29240 29404
rect 28976 29350 28986 29402
rect 29230 29350 29240 29402
rect 28976 29348 29000 29350
rect 29056 29348 29080 29350
rect 29136 29348 29160 29350
rect 29216 29348 29240 29350
rect 28920 29339 29296 29348
rect 22180 28860 22556 28869
rect 22236 28858 22260 28860
rect 22316 28858 22340 28860
rect 22396 28858 22420 28860
rect 22476 28858 22500 28860
rect 22236 28806 22246 28858
rect 22490 28806 22500 28858
rect 22236 28804 22260 28806
rect 22316 28804 22340 28806
rect 22396 28804 22420 28806
rect 22476 28804 22500 28806
rect 22180 28795 22556 28804
rect 28180 28860 28556 28869
rect 28236 28858 28260 28860
rect 28316 28858 28340 28860
rect 28396 28858 28420 28860
rect 28476 28858 28500 28860
rect 28236 28806 28246 28858
rect 28490 28806 28500 28858
rect 28236 28804 28260 28806
rect 28316 28804 28340 28806
rect 28396 28804 28420 28806
rect 28476 28804 28500 28806
rect 28180 28795 28556 28804
rect 22920 28316 23296 28325
rect 22976 28314 23000 28316
rect 23056 28314 23080 28316
rect 23136 28314 23160 28316
rect 23216 28314 23240 28316
rect 22976 28262 22986 28314
rect 23230 28262 23240 28314
rect 22976 28260 23000 28262
rect 23056 28260 23080 28262
rect 23136 28260 23160 28262
rect 23216 28260 23240 28262
rect 22920 28251 23296 28260
rect 28920 28316 29296 28325
rect 28976 28314 29000 28316
rect 29056 28314 29080 28316
rect 29136 28314 29160 28316
rect 29216 28314 29240 28316
rect 28976 28262 28986 28314
rect 29230 28262 29240 28314
rect 28976 28260 29000 28262
rect 29056 28260 29080 28262
rect 29136 28260 29160 28262
rect 29216 28260 29240 28262
rect 28920 28251 29296 28260
rect 23388 28076 23440 28082
rect 23388 28018 23440 28024
rect 26608 28076 26660 28082
rect 26608 28018 26660 28024
rect 20720 27940 20772 27946
rect 20720 27882 20772 27888
rect 20732 27470 20760 27882
rect 23112 27872 23164 27878
rect 23112 27814 23164 27820
rect 22180 27772 22556 27781
rect 22236 27770 22260 27772
rect 22316 27770 22340 27772
rect 22396 27770 22420 27772
rect 22476 27770 22500 27772
rect 22236 27718 22246 27770
rect 22490 27718 22500 27770
rect 22236 27716 22260 27718
rect 22316 27716 22340 27718
rect 22396 27716 22420 27718
rect 22476 27716 22500 27718
rect 22180 27707 22556 27716
rect 23124 27470 23152 27814
rect 20720 27464 20772 27470
rect 20720 27406 20772 27412
rect 22836 27464 22888 27470
rect 22836 27406 22888 27412
rect 23112 27464 23164 27470
rect 23112 27406 23164 27412
rect 21088 27328 21140 27334
rect 21088 27270 21140 27276
rect 21100 27130 21128 27270
rect 21088 27124 21140 27130
rect 21088 27066 21140 27072
rect 20536 26988 20588 26994
rect 20536 26930 20588 26936
rect 20444 26920 20496 26926
rect 20444 26862 20496 26868
rect 20364 24262 20484 24290
rect 20548 24274 20576 26930
rect 21180 26784 21232 26790
rect 21180 26726 21232 26732
rect 21192 26042 21220 26726
rect 22180 26684 22556 26693
rect 22236 26682 22260 26684
rect 22316 26682 22340 26684
rect 22396 26682 22420 26684
rect 22476 26682 22500 26684
rect 22236 26630 22246 26682
rect 22490 26630 22500 26682
rect 22236 26628 22260 26630
rect 22316 26628 22340 26630
rect 22396 26628 22420 26630
rect 22476 26628 22500 26630
rect 22180 26619 22556 26628
rect 21180 26036 21232 26042
rect 21180 25978 21232 25984
rect 22008 26036 22060 26042
rect 22008 25978 22060 25984
rect 21548 25152 21600 25158
rect 21548 25094 21600 25100
rect 20456 24206 20484 24262
rect 20536 24268 20588 24274
rect 20536 24210 20588 24216
rect 21180 24268 21232 24274
rect 21180 24210 21232 24216
rect 20352 24200 20404 24206
rect 20352 24142 20404 24148
rect 20444 24200 20496 24206
rect 20444 24142 20496 24148
rect 20364 23866 20392 24142
rect 20352 23860 20404 23866
rect 20352 23802 20404 23808
rect 20456 23798 20484 24142
rect 20720 24132 20772 24138
rect 20720 24074 20772 24080
rect 20732 23866 20760 24074
rect 20720 23860 20772 23866
rect 20720 23802 20772 23808
rect 20996 23860 21048 23866
rect 20996 23802 21048 23808
rect 20444 23792 20496 23798
rect 20444 23734 20496 23740
rect 20352 23724 20404 23730
rect 20352 23666 20404 23672
rect 20364 23186 20392 23666
rect 21008 23662 21036 23802
rect 21192 23730 21220 24210
rect 21560 24206 21588 25094
rect 21456 24200 21508 24206
rect 21456 24142 21508 24148
rect 21548 24200 21600 24206
rect 21600 24160 21680 24188
rect 21548 24142 21600 24148
rect 21180 23724 21232 23730
rect 21180 23666 21232 23672
rect 21468 23662 21496 24142
rect 21652 23662 21680 24160
rect 20996 23656 21048 23662
rect 20996 23598 21048 23604
rect 21456 23656 21508 23662
rect 21456 23598 21508 23604
rect 21640 23656 21692 23662
rect 21640 23598 21692 23604
rect 20352 23180 20404 23186
rect 20352 23122 20404 23128
rect 20628 22976 20680 22982
rect 20628 22918 20680 22924
rect 20640 22794 20668 22918
rect 20640 22778 20852 22794
rect 20640 22772 20864 22778
rect 20640 22766 20812 22772
rect 20812 22714 20864 22720
rect 20904 22636 20956 22642
rect 20904 22578 20956 22584
rect 20916 22386 20944 22578
rect 20732 22358 20944 22386
rect 20732 21962 20760 22358
rect 21008 22094 21036 23598
rect 21088 23588 21140 23594
rect 21088 23530 21140 23536
rect 21100 23118 21128 23530
rect 21548 23316 21600 23322
rect 21548 23258 21600 23264
rect 21088 23112 21140 23118
rect 21088 23054 21140 23060
rect 21560 23050 21588 23258
rect 21652 23186 21680 23598
rect 21640 23180 21692 23186
rect 21640 23122 21692 23128
rect 21272 23044 21324 23050
rect 21272 22986 21324 22992
rect 21548 23044 21600 23050
rect 21548 22986 21600 22992
rect 21284 22438 21312 22986
rect 21456 22568 21508 22574
rect 21456 22510 21508 22516
rect 21272 22432 21324 22438
rect 21272 22374 21324 22380
rect 21284 22166 21312 22374
rect 21468 22234 21496 22510
rect 21456 22228 21508 22234
rect 21456 22170 21508 22176
rect 21272 22160 21324 22166
rect 21272 22102 21324 22108
rect 20916 22066 21036 22094
rect 20720 21956 20772 21962
rect 20720 21898 20772 21904
rect 20732 21593 20760 21898
rect 20718 21584 20774 21593
rect 20718 21519 20774 21528
rect 20732 20777 20760 21519
rect 20718 20768 20774 20777
rect 20718 20703 20774 20712
rect 20444 19916 20496 19922
rect 20444 19858 20496 19864
rect 20260 18216 20312 18222
rect 20260 18158 20312 18164
rect 20352 18216 20404 18222
rect 20352 18158 20404 18164
rect 20076 18080 20128 18086
rect 20076 18022 20128 18028
rect 19984 17740 20036 17746
rect 19984 17682 20036 17688
rect 19340 17672 19392 17678
rect 19340 17614 19392 17620
rect 19524 17672 19576 17678
rect 19524 17614 19576 17620
rect 19800 17672 19852 17678
rect 19800 17614 19852 17620
rect 19340 17536 19392 17542
rect 19340 17478 19392 17484
rect 19352 17338 19380 17478
rect 19340 17332 19392 17338
rect 19340 17274 19392 17280
rect 19812 17270 19840 17614
rect 19800 17264 19852 17270
rect 19800 17206 19852 17212
rect 19892 17060 19944 17066
rect 19892 17002 19944 17008
rect 19156 16788 19208 16794
rect 19156 16730 19208 16736
rect 18972 16584 19024 16590
rect 18972 16526 19024 16532
rect 18972 15156 19024 15162
rect 18892 15116 18972 15144
rect 18972 15098 19024 15104
rect 19168 14482 19196 16730
rect 19708 15428 19760 15434
rect 19708 15370 19760 15376
rect 19156 14476 19208 14482
rect 19156 14418 19208 14424
rect 19720 14074 19748 15370
rect 19904 14482 19932 17002
rect 19892 14476 19944 14482
rect 19892 14418 19944 14424
rect 19708 14068 19760 14074
rect 19708 14010 19760 14016
rect 18604 14000 18656 14006
rect 18604 13942 18656 13948
rect 19720 13394 19748 14010
rect 19708 13388 19760 13394
rect 19708 13330 19760 13336
rect 19904 12434 19932 14418
rect 19996 14006 20024 17682
rect 20272 17066 20300 18158
rect 20364 17610 20392 18158
rect 20456 17678 20484 19858
rect 20720 19848 20772 19854
rect 20720 19790 20772 19796
rect 20732 18970 20760 19790
rect 20720 18964 20772 18970
rect 20720 18906 20772 18912
rect 20732 17678 20760 18906
rect 20812 18080 20864 18086
rect 20812 18022 20864 18028
rect 20444 17672 20496 17678
rect 20444 17614 20496 17620
rect 20720 17672 20772 17678
rect 20720 17614 20772 17620
rect 20352 17604 20404 17610
rect 20352 17546 20404 17552
rect 20352 17264 20404 17270
rect 20352 17206 20404 17212
rect 20260 17060 20312 17066
rect 20260 17002 20312 17008
rect 20076 15496 20128 15502
rect 20076 15438 20128 15444
rect 20088 14822 20116 15438
rect 20168 14884 20220 14890
rect 20168 14826 20220 14832
rect 20076 14816 20128 14822
rect 20076 14758 20128 14764
rect 20088 14006 20116 14758
rect 20180 14074 20208 14826
rect 20260 14816 20312 14822
rect 20260 14758 20312 14764
rect 20272 14618 20300 14758
rect 20260 14612 20312 14618
rect 20260 14554 20312 14560
rect 20168 14068 20220 14074
rect 20168 14010 20220 14016
rect 20260 14068 20312 14074
rect 20364 14056 20392 17206
rect 20824 14822 20852 18022
rect 20916 17678 20944 22066
rect 21180 19848 21232 19854
rect 21180 19790 21232 19796
rect 20996 19712 21048 19718
rect 20996 19654 21048 19660
rect 21008 19514 21036 19654
rect 20996 19508 21048 19514
rect 20996 19450 21048 19456
rect 21192 18970 21220 19790
rect 21456 19712 21508 19718
rect 21456 19654 21508 19660
rect 21180 18964 21232 18970
rect 21180 18906 21232 18912
rect 21468 18766 21496 19654
rect 21456 18760 21508 18766
rect 21456 18702 21508 18708
rect 21180 18284 21232 18290
rect 21180 18226 21232 18232
rect 21192 17882 21220 18226
rect 21272 18216 21324 18222
rect 21272 18158 21324 18164
rect 21284 17882 21312 18158
rect 21180 17876 21232 17882
rect 21180 17818 21232 17824
rect 21272 17876 21324 17882
rect 21272 17818 21324 17824
rect 21560 17678 21588 22986
rect 21652 22234 21680 23122
rect 21732 22976 21784 22982
rect 21732 22918 21784 22924
rect 21744 22642 21772 22918
rect 21732 22636 21784 22642
rect 21732 22578 21784 22584
rect 21640 22228 21692 22234
rect 21640 22170 21692 22176
rect 21744 22098 21772 22578
rect 21732 22092 21784 22098
rect 21732 22034 21784 22040
rect 22020 19922 22048 25978
rect 22848 25906 22876 27406
rect 22920 27228 23296 27237
rect 22976 27226 23000 27228
rect 23056 27226 23080 27228
rect 23136 27226 23160 27228
rect 23216 27226 23240 27228
rect 22976 27174 22986 27226
rect 23230 27174 23240 27226
rect 22976 27172 23000 27174
rect 23056 27172 23080 27174
rect 23136 27172 23160 27174
rect 23216 27172 23240 27174
rect 22920 27163 23296 27172
rect 23400 27130 23428 28018
rect 26332 27872 26384 27878
rect 26332 27814 26384 27820
rect 26344 27470 26372 27814
rect 25320 27464 25372 27470
rect 25320 27406 25372 27412
rect 26332 27464 26384 27470
rect 26332 27406 26384 27412
rect 24216 27328 24268 27334
rect 24216 27270 24268 27276
rect 24400 27328 24452 27334
rect 24400 27270 24452 27276
rect 23388 27124 23440 27130
rect 23388 27066 23440 27072
rect 23754 27024 23810 27033
rect 23754 26959 23756 26968
rect 23808 26959 23810 26968
rect 23756 26930 23808 26936
rect 23480 26376 23532 26382
rect 23480 26318 23532 26324
rect 23664 26376 23716 26382
rect 23664 26318 23716 26324
rect 23388 26240 23440 26246
rect 23388 26182 23440 26188
rect 22920 26140 23296 26149
rect 22976 26138 23000 26140
rect 23056 26138 23080 26140
rect 23136 26138 23160 26140
rect 23216 26138 23240 26140
rect 22976 26086 22986 26138
rect 23230 26086 23240 26138
rect 22976 26084 23000 26086
rect 23056 26084 23080 26086
rect 23136 26084 23160 26086
rect 23216 26084 23240 26086
rect 22920 26075 23296 26084
rect 23400 26024 23428 26182
rect 23216 25996 23428 26024
rect 23216 25906 23244 25996
rect 22836 25900 22888 25906
rect 22836 25842 22888 25848
rect 23204 25900 23256 25906
rect 23204 25842 23256 25848
rect 22652 25832 22704 25838
rect 22652 25774 22704 25780
rect 22180 25596 22556 25605
rect 22236 25594 22260 25596
rect 22316 25594 22340 25596
rect 22396 25594 22420 25596
rect 22476 25594 22500 25596
rect 22236 25542 22246 25594
rect 22490 25542 22500 25594
rect 22236 25540 22260 25542
rect 22316 25540 22340 25542
rect 22396 25540 22420 25542
rect 22476 25540 22500 25542
rect 22180 25531 22556 25540
rect 22664 25498 22692 25774
rect 23492 25498 23520 26318
rect 23676 25498 23704 26318
rect 24032 26240 24084 26246
rect 24032 26182 24084 26188
rect 24044 25838 24072 26182
rect 24032 25832 24084 25838
rect 24032 25774 24084 25780
rect 22652 25492 22704 25498
rect 22652 25434 22704 25440
rect 23480 25492 23532 25498
rect 23480 25434 23532 25440
rect 23664 25492 23716 25498
rect 23664 25434 23716 25440
rect 24032 25356 24084 25362
rect 24032 25298 24084 25304
rect 22920 25052 23296 25061
rect 22976 25050 23000 25052
rect 23056 25050 23080 25052
rect 23136 25050 23160 25052
rect 23216 25050 23240 25052
rect 22976 24998 22986 25050
rect 23230 24998 23240 25050
rect 22976 24996 23000 24998
rect 23056 24996 23080 24998
rect 23136 24996 23160 24998
rect 23216 24996 23240 24998
rect 22920 24987 23296 24996
rect 22180 24508 22556 24517
rect 22236 24506 22260 24508
rect 22316 24506 22340 24508
rect 22396 24506 22420 24508
rect 22476 24506 22500 24508
rect 22236 24454 22246 24506
rect 22490 24454 22500 24506
rect 22236 24452 22260 24454
rect 22316 24452 22340 24454
rect 22396 24452 22420 24454
rect 22476 24452 22500 24454
rect 22180 24443 22556 24452
rect 23388 24200 23440 24206
rect 23388 24142 23440 24148
rect 22920 23964 23296 23973
rect 22976 23962 23000 23964
rect 23056 23962 23080 23964
rect 23136 23962 23160 23964
rect 23216 23962 23240 23964
rect 22976 23910 22986 23962
rect 23230 23910 23240 23962
rect 22976 23908 23000 23910
rect 23056 23908 23080 23910
rect 23136 23908 23160 23910
rect 23216 23908 23240 23910
rect 22920 23899 23296 23908
rect 22180 23420 22556 23429
rect 22236 23418 22260 23420
rect 22316 23418 22340 23420
rect 22396 23418 22420 23420
rect 22476 23418 22500 23420
rect 22236 23366 22246 23418
rect 22490 23366 22500 23418
rect 22236 23364 22260 23366
rect 22316 23364 22340 23366
rect 22396 23364 22420 23366
rect 22476 23364 22500 23366
rect 22180 23355 22556 23364
rect 22560 23112 22612 23118
rect 22560 23054 22612 23060
rect 22284 23044 22336 23050
rect 22284 22986 22336 22992
rect 22296 22574 22324 22986
rect 22572 22642 22600 23054
rect 22652 23044 22704 23050
rect 22652 22986 22704 22992
rect 22744 23044 22796 23050
rect 22744 22986 22796 22992
rect 22664 22642 22692 22986
rect 22560 22636 22612 22642
rect 22560 22578 22612 22584
rect 22652 22636 22704 22642
rect 22652 22578 22704 22584
rect 22284 22568 22336 22574
rect 22284 22510 22336 22516
rect 22180 22332 22556 22341
rect 22236 22330 22260 22332
rect 22316 22330 22340 22332
rect 22396 22330 22420 22332
rect 22476 22330 22500 22332
rect 22236 22278 22246 22330
rect 22490 22278 22500 22330
rect 22236 22276 22260 22278
rect 22316 22276 22340 22278
rect 22396 22276 22420 22278
rect 22476 22276 22500 22278
rect 22180 22267 22556 22276
rect 22180 21244 22556 21253
rect 22236 21242 22260 21244
rect 22316 21242 22340 21244
rect 22396 21242 22420 21244
rect 22476 21242 22500 21244
rect 22236 21190 22246 21242
rect 22490 21190 22500 21242
rect 22236 21188 22260 21190
rect 22316 21188 22340 21190
rect 22396 21188 22420 21190
rect 22476 21188 22500 21190
rect 22180 21179 22556 21188
rect 22180 20156 22556 20165
rect 22236 20154 22260 20156
rect 22316 20154 22340 20156
rect 22396 20154 22420 20156
rect 22476 20154 22500 20156
rect 22236 20102 22246 20154
rect 22490 20102 22500 20154
rect 22236 20100 22260 20102
rect 22316 20100 22340 20102
rect 22396 20100 22420 20102
rect 22476 20100 22500 20102
rect 22180 20091 22556 20100
rect 22008 19916 22060 19922
rect 22008 19858 22060 19864
rect 22756 19786 22784 22986
rect 22920 22876 23296 22885
rect 22976 22874 23000 22876
rect 23056 22874 23080 22876
rect 23136 22874 23160 22876
rect 23216 22874 23240 22876
rect 22976 22822 22986 22874
rect 23230 22822 23240 22874
rect 22976 22820 23000 22822
rect 23056 22820 23080 22822
rect 23136 22820 23160 22822
rect 23216 22820 23240 22822
rect 22920 22811 23296 22820
rect 22836 22704 22888 22710
rect 22836 22646 22888 22652
rect 22848 22098 22876 22646
rect 22836 22092 22888 22098
rect 22836 22034 22888 22040
rect 22920 21788 23296 21797
rect 22976 21786 23000 21788
rect 23056 21786 23080 21788
rect 23136 21786 23160 21788
rect 23216 21786 23240 21788
rect 22976 21734 22986 21786
rect 23230 21734 23240 21786
rect 22976 21732 23000 21734
rect 23056 21732 23080 21734
rect 23136 21732 23160 21734
rect 23216 21732 23240 21734
rect 22920 21723 23296 21732
rect 22920 20700 23296 20709
rect 22976 20698 23000 20700
rect 23056 20698 23080 20700
rect 23136 20698 23160 20700
rect 23216 20698 23240 20700
rect 22976 20646 22986 20698
rect 23230 20646 23240 20698
rect 22976 20644 23000 20646
rect 23056 20644 23080 20646
rect 23136 20644 23160 20646
rect 23216 20644 23240 20646
rect 22920 20635 23296 20644
rect 22836 19848 22888 19854
rect 22836 19790 22888 19796
rect 22744 19780 22796 19786
rect 22744 19722 22796 19728
rect 21640 19712 21692 19718
rect 21640 19654 21692 19660
rect 21652 18834 21680 19654
rect 22100 19508 22152 19514
rect 22100 19450 22152 19456
rect 22112 18834 22140 19450
rect 22652 19372 22704 19378
rect 22652 19314 22704 19320
rect 22180 19068 22556 19077
rect 22236 19066 22260 19068
rect 22316 19066 22340 19068
rect 22396 19066 22420 19068
rect 22476 19066 22500 19068
rect 22236 19014 22246 19066
rect 22490 19014 22500 19066
rect 22236 19012 22260 19014
rect 22316 19012 22340 19014
rect 22396 19012 22420 19014
rect 22476 19012 22500 19014
rect 22180 19003 22556 19012
rect 22468 18896 22520 18902
rect 22664 18850 22692 19314
rect 22848 19174 22876 19790
rect 22920 19612 23296 19621
rect 22976 19610 23000 19612
rect 23056 19610 23080 19612
rect 23136 19610 23160 19612
rect 23216 19610 23240 19612
rect 22976 19558 22986 19610
rect 23230 19558 23240 19610
rect 22976 19556 23000 19558
rect 23056 19556 23080 19558
rect 23136 19556 23160 19558
rect 23216 19556 23240 19558
rect 22920 19547 23296 19556
rect 22836 19168 22888 19174
rect 22836 19110 22888 19116
rect 23020 19168 23072 19174
rect 23020 19110 23072 19116
rect 22520 18844 22692 18850
rect 22468 18838 22692 18844
rect 21640 18828 21692 18834
rect 21640 18770 21692 18776
rect 22100 18828 22152 18834
rect 22480 18822 22692 18838
rect 22100 18770 22152 18776
rect 21652 18408 21680 18770
rect 22848 18714 22876 19110
rect 23032 18834 23060 19110
rect 23400 18850 23428 24142
rect 23572 23656 23624 23662
rect 23572 23598 23624 23604
rect 23480 22976 23532 22982
rect 23480 22918 23532 22924
rect 23492 22778 23520 22918
rect 23480 22772 23532 22778
rect 23480 22714 23532 22720
rect 23480 21956 23532 21962
rect 23480 21898 23532 21904
rect 23492 21690 23520 21898
rect 23480 21684 23532 21690
rect 23480 21626 23532 21632
rect 23020 18828 23072 18834
rect 23020 18770 23072 18776
rect 23216 18822 23428 18850
rect 23216 18766 23244 18822
rect 23204 18760 23256 18766
rect 22848 18698 23060 18714
rect 23584 18714 23612 23598
rect 23664 23112 23716 23118
rect 23664 23054 23716 23060
rect 23676 22778 23704 23054
rect 23664 22772 23716 22778
rect 23664 22714 23716 22720
rect 23848 22704 23900 22710
rect 23848 22646 23900 22652
rect 23664 21888 23716 21894
rect 23664 21830 23716 21836
rect 23676 21554 23704 21830
rect 23860 21622 23888 22646
rect 24044 22166 24072 25298
rect 24228 24818 24256 27270
rect 24412 27130 24440 27270
rect 24400 27124 24452 27130
rect 24400 27066 24452 27072
rect 25332 26926 25360 27406
rect 26620 27130 26648 28018
rect 28180 27772 28556 27781
rect 28236 27770 28260 27772
rect 28316 27770 28340 27772
rect 28396 27770 28420 27772
rect 28476 27770 28500 27772
rect 28236 27718 28246 27770
rect 28490 27718 28500 27770
rect 28236 27716 28260 27718
rect 28316 27716 28340 27718
rect 28396 27716 28420 27718
rect 28476 27716 28500 27718
rect 28180 27707 28556 27716
rect 30576 27606 30604 32166
rect 29368 27600 29420 27606
rect 29368 27542 29420 27548
rect 30564 27600 30616 27606
rect 30564 27542 30616 27548
rect 27252 27328 27304 27334
rect 27252 27270 27304 27276
rect 27528 27328 27580 27334
rect 27528 27270 27580 27276
rect 26608 27124 26660 27130
rect 26608 27066 26660 27072
rect 25228 26920 25280 26926
rect 25228 26862 25280 26868
rect 25320 26920 25372 26926
rect 25320 26862 25372 26868
rect 24492 26444 24544 26450
rect 24492 26386 24544 26392
rect 24308 26376 24360 26382
rect 24308 26318 24360 26324
rect 24320 25770 24348 26318
rect 24400 26240 24452 26246
rect 24400 26182 24452 26188
rect 24308 25764 24360 25770
rect 24308 25706 24360 25712
rect 24320 24886 24348 25706
rect 24412 25294 24440 26182
rect 24504 25362 24532 26386
rect 24492 25356 24544 25362
rect 24492 25298 24544 25304
rect 25136 25356 25188 25362
rect 25136 25298 25188 25304
rect 24400 25288 24452 25294
rect 24400 25230 24452 25236
rect 24308 24880 24360 24886
rect 24308 24822 24360 24828
rect 24216 24812 24268 24818
rect 24216 24754 24268 24760
rect 24124 24744 24176 24750
rect 24124 24686 24176 24692
rect 24136 23322 24164 24686
rect 24308 24676 24360 24682
rect 24308 24618 24360 24624
rect 24320 23866 24348 24618
rect 24768 24608 24820 24614
rect 24768 24550 24820 24556
rect 24780 24274 24808 24550
rect 24768 24268 24820 24274
rect 24768 24210 24820 24216
rect 24308 23860 24360 23866
rect 24308 23802 24360 23808
rect 24124 23316 24176 23322
rect 24124 23258 24176 23264
rect 24032 22160 24084 22166
rect 24032 22102 24084 22108
rect 24136 21622 24164 23258
rect 24216 21888 24268 21894
rect 24216 21830 24268 21836
rect 24228 21622 24256 21830
rect 23848 21616 23900 21622
rect 23848 21558 23900 21564
rect 24124 21616 24176 21622
rect 24124 21558 24176 21564
rect 24216 21616 24268 21622
rect 24216 21558 24268 21564
rect 23664 21548 23716 21554
rect 23664 21490 23716 21496
rect 23860 21146 23888 21558
rect 24320 21554 24348 23802
rect 24860 23248 24912 23254
rect 24860 23190 24912 23196
rect 24768 23112 24820 23118
rect 24768 23054 24820 23060
rect 24780 22438 24808 23054
rect 24768 22432 24820 22438
rect 24768 22374 24820 22380
rect 24780 22094 24808 22374
rect 24872 22098 24900 23190
rect 25148 22386 25176 25298
rect 25240 22574 25268 26862
rect 25332 26450 25360 26862
rect 25320 26444 25372 26450
rect 25320 26386 25372 26392
rect 25332 25974 25360 26386
rect 26148 26308 26200 26314
rect 26148 26250 26200 26256
rect 25596 26036 25648 26042
rect 25596 25978 25648 25984
rect 25320 25968 25372 25974
rect 25320 25910 25372 25916
rect 25332 23186 25360 25910
rect 25608 25770 25636 25978
rect 25596 25764 25648 25770
rect 25596 25706 25648 25712
rect 25504 25696 25556 25702
rect 25504 25638 25556 25644
rect 25780 25696 25832 25702
rect 25780 25638 25832 25644
rect 26056 25696 26108 25702
rect 26056 25638 26108 25644
rect 25516 25158 25544 25638
rect 25792 25362 25820 25638
rect 26068 25498 26096 25638
rect 26056 25492 26108 25498
rect 26056 25434 26108 25440
rect 25780 25356 25832 25362
rect 25780 25298 25832 25304
rect 25504 25152 25556 25158
rect 25504 25094 25556 25100
rect 25792 24954 25820 25298
rect 26160 25158 26188 26250
rect 26884 26240 26936 26246
rect 26884 26182 26936 26188
rect 26896 25838 26924 26182
rect 26792 25832 26844 25838
rect 26792 25774 26844 25780
rect 26884 25832 26936 25838
rect 26884 25774 26936 25780
rect 26804 25702 26832 25774
rect 26792 25696 26844 25702
rect 26792 25638 26844 25644
rect 26148 25152 26200 25158
rect 26148 25094 26200 25100
rect 25780 24948 25832 24954
rect 25780 24890 25832 24896
rect 26516 24812 26568 24818
rect 26516 24754 26568 24760
rect 25964 24608 26016 24614
rect 25964 24550 26016 24556
rect 25976 24410 26004 24550
rect 25964 24404 26016 24410
rect 25964 24346 26016 24352
rect 26056 24200 26108 24206
rect 26056 24142 26108 24148
rect 26068 23866 26096 24142
rect 26528 24070 26556 24754
rect 26700 24676 26752 24682
rect 26700 24618 26752 24624
rect 26516 24064 26568 24070
rect 26516 24006 26568 24012
rect 26056 23860 26108 23866
rect 26056 23802 26108 23808
rect 26424 23724 26476 23730
rect 26424 23666 26476 23672
rect 26240 23520 26292 23526
rect 26240 23462 26292 23468
rect 25320 23180 25372 23186
rect 25320 23122 25372 23128
rect 26056 23112 26108 23118
rect 26056 23054 26108 23060
rect 25412 22976 25464 22982
rect 25412 22918 25464 22924
rect 25424 22778 25452 22918
rect 25412 22772 25464 22778
rect 25412 22714 25464 22720
rect 25228 22568 25280 22574
rect 25228 22510 25280 22516
rect 25148 22358 25268 22386
rect 24688 22066 24808 22094
rect 24860 22092 24912 22098
rect 24308 21548 24360 21554
rect 24308 21490 24360 21496
rect 24688 21486 24716 22066
rect 24912 22052 24992 22080
rect 24860 22034 24912 22040
rect 24768 21888 24820 21894
rect 24768 21830 24820 21836
rect 24780 21690 24808 21830
rect 24768 21684 24820 21690
rect 24768 21626 24820 21632
rect 24860 21616 24912 21622
rect 24858 21584 24860 21593
rect 24912 21584 24914 21593
rect 24858 21519 24914 21528
rect 24676 21480 24728 21486
rect 24676 21422 24728 21428
rect 23848 21140 23900 21146
rect 23848 21082 23900 21088
rect 24964 21010 24992 22052
rect 24952 21004 25004 21010
rect 24952 20946 25004 20952
rect 24964 20466 24992 20946
rect 25044 20936 25096 20942
rect 25044 20878 25096 20884
rect 25056 20602 25084 20878
rect 25044 20596 25096 20602
rect 25044 20538 25096 20544
rect 23940 20460 23992 20466
rect 23940 20402 23992 20408
rect 24952 20460 25004 20466
rect 24952 20402 25004 20408
rect 23952 20058 23980 20402
rect 25240 20398 25268 22358
rect 25320 21956 25372 21962
rect 25320 21898 25372 21904
rect 25332 21622 25360 21898
rect 26068 21622 26096 23054
rect 26252 23050 26280 23462
rect 26240 23044 26292 23050
rect 26240 22986 26292 22992
rect 26436 22098 26464 23666
rect 26424 22092 26476 22098
rect 26424 22034 26476 22040
rect 26148 21956 26200 21962
rect 26148 21898 26200 21904
rect 25320 21616 25372 21622
rect 25320 21558 25372 21564
rect 26056 21616 26108 21622
rect 26056 21558 26108 21564
rect 25320 20800 25372 20806
rect 25320 20742 25372 20748
rect 25332 20602 25360 20742
rect 25320 20596 25372 20602
rect 25320 20538 25372 20544
rect 26160 20534 26188 21898
rect 26240 21888 26292 21894
rect 26240 21830 26292 21836
rect 26148 20528 26200 20534
rect 26148 20470 26200 20476
rect 25228 20392 25280 20398
rect 25228 20334 25280 20340
rect 25136 20256 25188 20262
rect 25136 20198 25188 20204
rect 25148 20058 25176 20198
rect 23940 20052 23992 20058
rect 23940 19994 23992 20000
rect 25136 20052 25188 20058
rect 25136 19994 25188 20000
rect 23664 19780 23716 19786
rect 23664 19722 23716 19728
rect 23204 18702 23256 18708
rect 23400 18698 23612 18714
rect 22848 18692 23072 18698
rect 22848 18686 23020 18692
rect 23020 18634 23072 18640
rect 23388 18692 23612 18698
rect 23440 18686 23612 18692
rect 23388 18634 23440 18640
rect 22744 18624 22796 18630
rect 22744 18566 22796 18572
rect 22836 18624 22888 18630
rect 22836 18566 22888 18572
rect 21732 18420 21784 18426
rect 21652 18380 21732 18408
rect 21652 18154 21680 18380
rect 21732 18362 21784 18368
rect 22756 18222 22784 18566
rect 22744 18216 22796 18222
rect 22744 18158 22796 18164
rect 21640 18148 21692 18154
rect 21640 18090 21692 18096
rect 22180 17980 22556 17989
rect 22236 17978 22260 17980
rect 22316 17978 22340 17980
rect 22396 17978 22420 17980
rect 22476 17978 22500 17980
rect 22236 17926 22246 17978
rect 22490 17926 22500 17978
rect 22236 17924 22260 17926
rect 22316 17924 22340 17926
rect 22396 17924 22420 17926
rect 22476 17924 22500 17926
rect 22180 17915 22556 17924
rect 20904 17672 20956 17678
rect 20904 17614 20956 17620
rect 21548 17672 21600 17678
rect 21548 17614 21600 17620
rect 20916 15502 20944 17614
rect 21732 17604 21784 17610
rect 21732 17546 21784 17552
rect 21548 16584 21600 16590
rect 21548 16526 21600 16532
rect 21560 16046 21588 16526
rect 21744 16250 21772 17546
rect 22652 17196 22704 17202
rect 22652 17138 22704 17144
rect 22100 16992 22152 16998
rect 22100 16934 22152 16940
rect 22112 16590 22140 16934
rect 22180 16892 22556 16901
rect 22236 16890 22260 16892
rect 22316 16890 22340 16892
rect 22396 16890 22420 16892
rect 22476 16890 22500 16892
rect 22236 16838 22246 16890
rect 22490 16838 22500 16890
rect 22236 16836 22260 16838
rect 22316 16836 22340 16838
rect 22396 16836 22420 16838
rect 22476 16836 22500 16838
rect 22180 16827 22556 16836
rect 22100 16584 22152 16590
rect 22100 16526 22152 16532
rect 21732 16244 21784 16250
rect 21732 16186 21784 16192
rect 21364 16040 21416 16046
rect 21362 16008 21364 16017
rect 21548 16040 21600 16046
rect 21416 16008 21418 16017
rect 21548 15982 21600 15988
rect 21362 15943 21418 15952
rect 21180 15904 21232 15910
rect 21180 15846 21232 15852
rect 20904 15496 20956 15502
rect 20904 15438 20956 15444
rect 20996 15496 21048 15502
rect 20996 15438 21048 15444
rect 20904 15360 20956 15366
rect 20904 15302 20956 15308
rect 20812 14816 20864 14822
rect 20812 14758 20864 14764
rect 20312 14028 20392 14056
rect 20260 14010 20312 14016
rect 19984 14000 20036 14006
rect 19984 13942 20036 13948
rect 20076 14000 20128 14006
rect 20076 13942 20128 13948
rect 19812 12406 19932 12434
rect 19248 12096 19300 12102
rect 19248 12038 19300 12044
rect 19708 12096 19760 12102
rect 19708 12038 19760 12044
rect 18972 11552 19024 11558
rect 18972 11494 19024 11500
rect 18984 9586 19012 11494
rect 19260 11150 19288 12038
rect 19432 11756 19484 11762
rect 19432 11698 19484 11704
rect 19444 11354 19472 11698
rect 19432 11348 19484 11354
rect 19432 11290 19484 11296
rect 19248 11144 19300 11150
rect 19248 11086 19300 11092
rect 19720 11014 19748 12038
rect 19432 11008 19484 11014
rect 19432 10950 19484 10956
rect 19708 11008 19760 11014
rect 19708 10950 19760 10956
rect 19444 9926 19472 10950
rect 19524 10668 19576 10674
rect 19524 10610 19576 10616
rect 19340 9920 19392 9926
rect 19340 9862 19392 9868
rect 19432 9920 19484 9926
rect 19432 9862 19484 9868
rect 18972 9580 19024 9586
rect 18972 9522 19024 9528
rect 18512 9172 18564 9178
rect 18512 9114 18564 9120
rect 18984 8974 19012 9522
rect 19248 9376 19300 9382
rect 19352 9330 19380 9862
rect 19444 9586 19472 9862
rect 19432 9580 19484 9586
rect 19432 9522 19484 9528
rect 19300 9324 19380 9330
rect 19248 9318 19380 9324
rect 19260 9302 19380 9318
rect 19444 9194 19472 9522
rect 19168 9166 19472 9194
rect 18512 8968 18564 8974
rect 18512 8910 18564 8916
rect 18972 8968 19024 8974
rect 18972 8910 19024 8916
rect 18052 8900 18104 8906
rect 18052 8842 18104 8848
rect 18064 8634 18092 8842
rect 18052 8628 18104 8634
rect 18052 8570 18104 8576
rect 18524 8362 18552 8910
rect 18696 8900 18748 8906
rect 18696 8842 18748 8848
rect 18708 8566 18736 8842
rect 19168 8634 19196 9166
rect 19340 9104 19392 9110
rect 19340 9046 19392 9052
rect 19156 8628 19208 8634
rect 19156 8570 19208 8576
rect 18696 8560 18748 8566
rect 18696 8502 18748 8508
rect 18512 8356 18564 8362
rect 18512 8298 18564 8304
rect 18524 8090 18552 8298
rect 19352 8090 19380 9046
rect 19432 8900 19484 8906
rect 19432 8842 19484 8848
rect 19444 8634 19472 8842
rect 19432 8628 19484 8634
rect 19432 8570 19484 8576
rect 19432 8424 19484 8430
rect 19432 8366 19484 8372
rect 18512 8084 18564 8090
rect 18512 8026 18564 8032
rect 19340 8084 19392 8090
rect 19340 8026 19392 8032
rect 19444 8022 19472 8366
rect 19432 8016 19484 8022
rect 19432 7958 19484 7964
rect 19432 6928 19484 6934
rect 19432 6870 19484 6876
rect 19156 6792 19208 6798
rect 19156 6734 19208 6740
rect 18788 6656 18840 6662
rect 18788 6598 18840 6604
rect 19064 6656 19116 6662
rect 19064 6598 19116 6604
rect 16764 6248 16816 6254
rect 16764 6190 16816 6196
rect 17868 6248 17920 6254
rect 17868 6190 17920 6196
rect 17408 6112 17460 6118
rect 17408 6054 17460 6060
rect 16672 5772 16724 5778
rect 16672 5714 16724 5720
rect 17316 5636 17368 5642
rect 17316 5578 17368 5584
rect 16920 5468 17296 5477
rect 16976 5466 17000 5468
rect 17056 5466 17080 5468
rect 17136 5466 17160 5468
rect 17216 5466 17240 5468
rect 16976 5414 16986 5466
rect 17230 5414 17240 5466
rect 16976 5412 17000 5414
rect 17056 5412 17080 5414
rect 17136 5412 17160 5414
rect 17216 5412 17240 5414
rect 16920 5403 17296 5412
rect 17328 5370 17356 5578
rect 17420 5370 17448 6054
rect 17880 5778 17908 6190
rect 18236 6112 18288 6118
rect 18236 6054 18288 6060
rect 18248 5914 18276 6054
rect 18236 5908 18288 5914
rect 18236 5850 18288 5856
rect 18800 5778 18828 6598
rect 19076 6390 19104 6598
rect 19168 6458 19196 6734
rect 19156 6452 19208 6458
rect 19156 6394 19208 6400
rect 19064 6384 19116 6390
rect 19064 6326 19116 6332
rect 19248 6384 19300 6390
rect 19444 6338 19472 6870
rect 19536 6458 19564 10610
rect 19708 10600 19760 10606
rect 19708 10542 19760 10548
rect 19720 9178 19748 10542
rect 19708 9172 19760 9178
rect 19708 9114 19760 9120
rect 19812 8022 19840 12406
rect 19892 8968 19944 8974
rect 19892 8910 19944 8916
rect 19800 8016 19852 8022
rect 19800 7958 19852 7964
rect 19616 7744 19668 7750
rect 19616 7686 19668 7692
rect 19628 7546 19656 7686
rect 19616 7540 19668 7546
rect 19616 7482 19668 7488
rect 19904 7478 19932 8910
rect 19996 8566 20024 13942
rect 20364 12434 20392 14028
rect 20824 13870 20852 14758
rect 20916 14618 20944 15302
rect 21008 14958 21036 15438
rect 21192 15366 21220 15846
rect 21180 15360 21232 15366
rect 21180 15302 21232 15308
rect 21560 15094 21588 15982
rect 21744 15638 21772 16186
rect 22100 15904 22152 15910
rect 22100 15846 22152 15852
rect 21732 15632 21784 15638
rect 21784 15580 22048 15586
rect 21732 15574 22048 15580
rect 21744 15558 22048 15574
rect 21548 15088 21600 15094
rect 21548 15030 21600 15036
rect 21272 15020 21324 15026
rect 21272 14962 21324 14968
rect 20996 14952 21048 14958
rect 20996 14894 21048 14900
rect 20904 14612 20956 14618
rect 20904 14554 20956 14560
rect 21008 14278 21036 14894
rect 20996 14272 21048 14278
rect 20996 14214 21048 14220
rect 21088 14272 21140 14278
rect 21088 14214 21140 14220
rect 21100 13938 21128 14214
rect 21088 13932 21140 13938
rect 21088 13874 21140 13880
rect 21284 13870 21312 14962
rect 21364 14884 21416 14890
rect 21364 14826 21416 14832
rect 21376 14414 21404 14826
rect 21560 14414 21588 15030
rect 21640 14816 21692 14822
rect 21640 14758 21692 14764
rect 21364 14408 21416 14414
rect 21548 14408 21600 14414
rect 21364 14350 21416 14356
rect 21468 14356 21548 14362
rect 21468 14350 21600 14356
rect 21468 14334 21588 14350
rect 20812 13864 20864 13870
rect 20812 13806 20864 13812
rect 21272 13864 21324 13870
rect 21272 13806 21324 13812
rect 20536 12844 20588 12850
rect 20536 12786 20588 12792
rect 20442 12744 20498 12753
rect 20548 12730 20576 12786
rect 21468 12782 21496 14334
rect 21652 14074 21680 14758
rect 21732 14612 21784 14618
rect 21732 14554 21784 14560
rect 21640 14068 21692 14074
rect 21640 14010 21692 14016
rect 21744 13938 21772 14554
rect 21732 13932 21784 13938
rect 21732 13874 21784 13880
rect 21732 13728 21784 13734
rect 21732 13670 21784 13676
rect 20498 12702 20576 12730
rect 21456 12776 21508 12782
rect 21456 12718 21508 12724
rect 20442 12679 20498 12688
rect 20548 12434 20576 12702
rect 20364 12406 20484 12434
rect 20548 12406 20760 12434
rect 20352 11552 20404 11558
rect 20352 11494 20404 11500
rect 20364 11218 20392 11494
rect 20352 11212 20404 11218
rect 20352 11154 20404 11160
rect 20260 10668 20312 10674
rect 20260 10610 20312 10616
rect 20352 10668 20404 10674
rect 20352 10610 20404 10616
rect 20076 10464 20128 10470
rect 20076 10406 20128 10412
rect 20168 10464 20220 10470
rect 20168 10406 20220 10412
rect 20088 10266 20116 10406
rect 20076 10260 20128 10266
rect 20076 10202 20128 10208
rect 20180 8974 20208 10406
rect 20272 10266 20300 10610
rect 20260 10260 20312 10266
rect 20260 10202 20312 10208
rect 20260 10056 20312 10062
rect 20260 9998 20312 10004
rect 20272 9722 20300 9998
rect 20364 9722 20392 10610
rect 20260 9716 20312 9722
rect 20260 9658 20312 9664
rect 20352 9716 20404 9722
rect 20352 9658 20404 9664
rect 20168 8968 20220 8974
rect 20168 8910 20220 8916
rect 20456 8634 20484 12406
rect 20732 11830 20760 12406
rect 21468 12306 21496 12718
rect 21744 12434 21772 13670
rect 21744 12406 21956 12434
rect 21456 12300 21508 12306
rect 21456 12242 21508 12248
rect 21272 12164 21324 12170
rect 21272 12106 21324 12112
rect 21088 12096 21140 12102
rect 21088 12038 21140 12044
rect 20720 11824 20772 11830
rect 20720 11766 20772 11772
rect 21100 11558 21128 12038
rect 21088 11552 21140 11558
rect 21088 11494 21140 11500
rect 21180 11552 21232 11558
rect 21180 11494 21232 11500
rect 21100 11082 21128 11494
rect 21192 11082 21220 11494
rect 21284 11354 21312 12106
rect 21640 11824 21692 11830
rect 21638 11792 21640 11801
rect 21692 11792 21694 11801
rect 21638 11727 21694 11736
rect 21272 11348 21324 11354
rect 21272 11290 21324 11296
rect 21088 11076 21140 11082
rect 21088 11018 21140 11024
rect 21180 11076 21232 11082
rect 21180 11018 21232 11024
rect 20812 11008 20864 11014
rect 20812 10950 20864 10956
rect 20824 10470 20852 10950
rect 20812 10464 20864 10470
rect 20812 10406 20864 10412
rect 21180 9988 21232 9994
rect 21180 9930 21232 9936
rect 21272 9988 21324 9994
rect 21272 9930 21324 9936
rect 20720 9580 20772 9586
rect 20720 9522 20772 9528
rect 20732 9178 20760 9522
rect 20720 9172 20772 9178
rect 20720 9114 20772 9120
rect 21192 9042 21220 9930
rect 21284 9722 21312 9930
rect 21272 9716 21324 9722
rect 21272 9658 21324 9664
rect 21180 9036 21232 9042
rect 21180 8978 21232 8984
rect 21824 9036 21876 9042
rect 21824 8978 21876 8984
rect 20444 8628 20496 8634
rect 20444 8570 20496 8576
rect 19984 8560 20036 8566
rect 19984 8502 20036 8508
rect 21836 8294 21864 8978
rect 21744 8266 21864 8294
rect 20628 8084 20680 8090
rect 20628 8026 20680 8032
rect 20640 7954 20668 8026
rect 20628 7948 20680 7954
rect 20628 7890 20680 7896
rect 20628 7744 20680 7750
rect 20628 7686 20680 7692
rect 21640 7744 21692 7750
rect 21640 7686 21692 7692
rect 19892 7472 19944 7478
rect 19892 7414 19944 7420
rect 19524 6452 19576 6458
rect 19524 6394 19576 6400
rect 19708 6452 19760 6458
rect 19708 6394 19760 6400
rect 19248 6326 19300 6332
rect 19260 5778 19288 6326
rect 19398 6322 19472 6338
rect 19386 6316 19472 6322
rect 19438 6310 19472 6316
rect 19386 6258 19438 6264
rect 17868 5772 17920 5778
rect 17868 5714 17920 5720
rect 18788 5772 18840 5778
rect 18788 5714 18840 5720
rect 19248 5772 19300 5778
rect 19248 5714 19300 5720
rect 18880 5704 18932 5710
rect 18880 5646 18932 5652
rect 18328 5568 18380 5574
rect 18328 5510 18380 5516
rect 17316 5364 17368 5370
rect 17316 5306 17368 5312
rect 17408 5364 17460 5370
rect 17408 5306 17460 5312
rect 17776 5228 17828 5234
rect 17776 5170 17828 5176
rect 16180 4924 16556 4933
rect 16236 4922 16260 4924
rect 16316 4922 16340 4924
rect 16396 4922 16420 4924
rect 16476 4922 16500 4924
rect 16236 4870 16246 4922
rect 16490 4870 16500 4922
rect 16236 4868 16260 4870
rect 16316 4868 16340 4870
rect 16396 4868 16420 4870
rect 16476 4868 16500 4870
rect 16180 4859 16556 4868
rect 17788 4826 17816 5170
rect 17776 4820 17828 4826
rect 17776 4762 17828 4768
rect 18340 4622 18368 5510
rect 18892 5370 18920 5646
rect 19720 5574 19748 6394
rect 19708 5568 19760 5574
rect 19708 5510 19760 5516
rect 19800 5568 19852 5574
rect 19800 5510 19852 5516
rect 18880 5364 18932 5370
rect 18880 5306 18932 5312
rect 19812 5234 19840 5510
rect 19904 5234 19932 7414
rect 20640 6730 20668 7686
rect 21652 7410 21680 7686
rect 21640 7404 21692 7410
rect 21640 7346 21692 7352
rect 21744 6934 21772 8266
rect 21824 7880 21876 7886
rect 21824 7822 21876 7828
rect 21732 6928 21784 6934
rect 21732 6870 21784 6876
rect 20812 6860 20864 6866
rect 20812 6802 20864 6808
rect 20628 6724 20680 6730
rect 20628 6666 20680 6672
rect 20640 5778 20668 6666
rect 20824 5778 20852 6802
rect 21836 6662 21864 7822
rect 21824 6656 21876 6662
rect 21824 6598 21876 6604
rect 21548 6248 21600 6254
rect 21548 6190 21600 6196
rect 20996 6112 21048 6118
rect 20996 6054 21048 6060
rect 21008 5914 21036 6054
rect 20996 5908 21048 5914
rect 20996 5850 21048 5856
rect 20628 5772 20680 5778
rect 20628 5714 20680 5720
rect 20812 5772 20864 5778
rect 20812 5714 20864 5720
rect 21272 5568 21324 5574
rect 21272 5510 21324 5516
rect 21284 5370 21312 5510
rect 21272 5364 21324 5370
rect 21272 5306 21324 5312
rect 19800 5228 19852 5234
rect 19800 5170 19852 5176
rect 19892 5228 19944 5234
rect 19892 5170 19944 5176
rect 19904 4690 19932 5170
rect 21560 5098 21588 6190
rect 21836 5914 21864 6598
rect 21824 5908 21876 5914
rect 21824 5850 21876 5856
rect 21928 5794 21956 12406
rect 22020 6730 22048 15558
rect 22112 15162 22140 15846
rect 22180 15804 22556 15813
rect 22236 15802 22260 15804
rect 22316 15802 22340 15804
rect 22396 15802 22420 15804
rect 22476 15802 22500 15804
rect 22236 15750 22246 15802
rect 22490 15750 22500 15802
rect 22236 15748 22260 15750
rect 22316 15748 22340 15750
rect 22396 15748 22420 15750
rect 22476 15748 22500 15750
rect 22180 15739 22556 15748
rect 22664 15706 22692 17138
rect 22744 16992 22796 16998
rect 22744 16934 22796 16940
rect 22376 15700 22428 15706
rect 22376 15642 22428 15648
rect 22652 15700 22704 15706
rect 22652 15642 22704 15648
rect 22100 15156 22152 15162
rect 22100 15098 22152 15104
rect 22388 15026 22416 15642
rect 22560 15632 22612 15638
rect 22480 15592 22560 15620
rect 22480 15502 22508 15592
rect 22560 15574 22612 15580
rect 22468 15496 22520 15502
rect 22468 15438 22520 15444
rect 22480 15042 22508 15438
rect 22756 15162 22784 16934
rect 22744 15156 22796 15162
rect 22744 15098 22796 15104
rect 22376 15020 22428 15026
rect 22480 15014 22784 15042
rect 22376 14962 22428 14968
rect 22180 14716 22556 14725
rect 22236 14714 22260 14716
rect 22316 14714 22340 14716
rect 22396 14714 22420 14716
rect 22476 14714 22500 14716
rect 22236 14662 22246 14714
rect 22490 14662 22500 14714
rect 22236 14660 22260 14662
rect 22316 14660 22340 14662
rect 22396 14660 22420 14662
rect 22476 14660 22500 14662
rect 22180 14651 22556 14660
rect 22100 14068 22152 14074
rect 22100 14010 22152 14016
rect 22112 13462 22140 14010
rect 22652 13796 22704 13802
rect 22652 13738 22704 13744
rect 22180 13628 22556 13637
rect 22236 13626 22260 13628
rect 22316 13626 22340 13628
rect 22396 13626 22420 13628
rect 22476 13626 22500 13628
rect 22236 13574 22246 13626
rect 22490 13574 22500 13626
rect 22236 13572 22260 13574
rect 22316 13572 22340 13574
rect 22396 13572 22420 13574
rect 22476 13572 22500 13574
rect 22180 13563 22556 13572
rect 22100 13456 22152 13462
rect 22100 13398 22152 13404
rect 22664 12986 22692 13738
rect 22652 12980 22704 12986
rect 22652 12922 22704 12928
rect 22100 12640 22152 12646
rect 22100 12582 22152 12588
rect 22112 11830 22140 12582
rect 22180 12540 22556 12549
rect 22236 12538 22260 12540
rect 22316 12538 22340 12540
rect 22396 12538 22420 12540
rect 22476 12538 22500 12540
rect 22236 12486 22246 12538
rect 22490 12486 22500 12538
rect 22236 12484 22260 12486
rect 22316 12484 22340 12486
rect 22396 12484 22420 12486
rect 22476 12484 22500 12486
rect 22180 12475 22556 12484
rect 22756 12434 22784 15014
rect 22664 12406 22784 12434
rect 22100 11824 22152 11830
rect 22100 11766 22152 11772
rect 22284 11824 22336 11830
rect 22284 11766 22336 11772
rect 22296 11642 22324 11766
rect 22112 11614 22324 11642
rect 22112 11218 22140 11614
rect 22180 11452 22556 11461
rect 22236 11450 22260 11452
rect 22316 11450 22340 11452
rect 22396 11450 22420 11452
rect 22476 11450 22500 11452
rect 22236 11398 22246 11450
rect 22490 11398 22500 11450
rect 22236 11396 22260 11398
rect 22316 11396 22340 11398
rect 22396 11396 22420 11398
rect 22476 11396 22500 11398
rect 22180 11387 22556 11396
rect 22100 11212 22152 11218
rect 22100 11154 22152 11160
rect 22180 10364 22556 10373
rect 22236 10362 22260 10364
rect 22316 10362 22340 10364
rect 22396 10362 22420 10364
rect 22476 10362 22500 10364
rect 22236 10310 22246 10362
rect 22490 10310 22500 10362
rect 22236 10308 22260 10310
rect 22316 10308 22340 10310
rect 22396 10308 22420 10310
rect 22476 10308 22500 10310
rect 22180 10299 22556 10308
rect 22180 9276 22556 9285
rect 22236 9274 22260 9276
rect 22316 9274 22340 9276
rect 22396 9274 22420 9276
rect 22476 9274 22500 9276
rect 22236 9222 22246 9274
rect 22490 9222 22500 9274
rect 22236 9220 22260 9222
rect 22316 9220 22340 9222
rect 22396 9220 22420 9222
rect 22476 9220 22500 9222
rect 22180 9211 22556 9220
rect 22664 9042 22692 12406
rect 22848 12186 22876 18566
rect 22920 18524 23296 18533
rect 22976 18522 23000 18524
rect 23056 18522 23080 18524
rect 23136 18522 23160 18524
rect 23216 18522 23240 18524
rect 22976 18470 22986 18522
rect 23230 18470 23240 18522
rect 22976 18468 23000 18470
rect 23056 18468 23080 18470
rect 23136 18468 23160 18470
rect 23216 18468 23240 18470
rect 22920 18459 23296 18468
rect 22920 17436 23296 17445
rect 22976 17434 23000 17436
rect 23056 17434 23080 17436
rect 23136 17434 23160 17436
rect 23216 17434 23240 17436
rect 22976 17382 22986 17434
rect 23230 17382 23240 17434
rect 22976 17380 23000 17382
rect 23056 17380 23080 17382
rect 23136 17380 23160 17382
rect 23216 17380 23240 17382
rect 22920 17371 23296 17380
rect 23400 16538 23428 18634
rect 23572 17128 23624 17134
rect 23572 17070 23624 17076
rect 23400 16510 23520 16538
rect 23388 16448 23440 16454
rect 23388 16390 23440 16396
rect 22920 16348 23296 16357
rect 22976 16346 23000 16348
rect 23056 16346 23080 16348
rect 23136 16346 23160 16348
rect 23216 16346 23240 16348
rect 22976 16294 22986 16346
rect 23230 16294 23240 16346
rect 22976 16292 23000 16294
rect 23056 16292 23080 16294
rect 23136 16292 23160 16294
rect 23216 16292 23240 16294
rect 22920 16283 23296 16292
rect 23400 16182 23428 16390
rect 23388 16176 23440 16182
rect 23388 16118 23440 16124
rect 23204 16108 23256 16114
rect 23204 16050 23256 16056
rect 22926 16008 22982 16017
rect 22926 15943 22982 15952
rect 22940 15570 22968 15943
rect 23216 15638 23244 16050
rect 23400 15706 23428 16118
rect 23388 15700 23440 15706
rect 23388 15642 23440 15648
rect 23204 15632 23256 15638
rect 23492 15586 23520 16510
rect 23584 16182 23612 17070
rect 23572 16176 23624 16182
rect 23572 16118 23624 16124
rect 23584 15978 23612 16118
rect 23572 15972 23624 15978
rect 23572 15914 23624 15920
rect 23204 15574 23256 15580
rect 22928 15564 22980 15570
rect 22928 15506 22980 15512
rect 23020 15564 23072 15570
rect 23020 15506 23072 15512
rect 23400 15558 23520 15586
rect 23032 15366 23060 15506
rect 23020 15360 23072 15366
rect 23020 15302 23072 15308
rect 22920 15260 23296 15269
rect 22976 15258 23000 15260
rect 23056 15258 23080 15260
rect 23136 15258 23160 15260
rect 23216 15258 23240 15260
rect 22976 15206 22986 15258
rect 23230 15206 23240 15258
rect 22976 15204 23000 15206
rect 23056 15204 23080 15206
rect 23136 15204 23160 15206
rect 23216 15204 23240 15206
rect 22920 15195 23296 15204
rect 22920 14172 23296 14181
rect 22976 14170 23000 14172
rect 23056 14170 23080 14172
rect 23136 14170 23160 14172
rect 23216 14170 23240 14172
rect 22976 14118 22986 14170
rect 23230 14118 23240 14170
rect 22976 14116 23000 14118
rect 23056 14116 23080 14118
rect 23136 14116 23160 14118
rect 23216 14116 23240 14118
rect 22920 14107 23296 14116
rect 23296 13932 23348 13938
rect 23296 13874 23348 13880
rect 23308 13530 23336 13874
rect 23296 13524 23348 13530
rect 23296 13466 23348 13472
rect 22920 13084 23296 13093
rect 22976 13082 23000 13084
rect 23056 13082 23080 13084
rect 23136 13082 23160 13084
rect 23216 13082 23240 13084
rect 22976 13030 22986 13082
rect 23230 13030 23240 13082
rect 22976 13028 23000 13030
rect 23056 13028 23080 13030
rect 23136 13028 23160 13030
rect 23216 13028 23240 13030
rect 22920 13019 23296 13028
rect 22928 12844 22980 12850
rect 22928 12786 22980 12792
rect 22940 12442 22968 12786
rect 23296 12640 23348 12646
rect 23296 12582 23348 12588
rect 22928 12436 22980 12442
rect 22928 12378 22980 12384
rect 23308 12238 23336 12582
rect 22756 12158 22876 12186
rect 23296 12232 23348 12238
rect 23296 12174 23348 12180
rect 22756 11150 22784 12158
rect 22836 12096 22888 12102
rect 22836 12038 22888 12044
rect 22848 11762 22876 12038
rect 22920 11996 23296 12005
rect 22976 11994 23000 11996
rect 23056 11994 23080 11996
rect 23136 11994 23160 11996
rect 23216 11994 23240 11996
rect 22976 11942 22986 11994
rect 23230 11942 23240 11994
rect 22976 11940 23000 11942
rect 23056 11940 23080 11942
rect 23136 11940 23160 11942
rect 23216 11940 23240 11942
rect 22920 11931 23296 11940
rect 22836 11756 22888 11762
rect 22836 11698 22888 11704
rect 23400 11558 23428 15558
rect 23480 11756 23532 11762
rect 23480 11698 23532 11704
rect 23388 11552 23440 11558
rect 23388 11494 23440 11500
rect 22836 11348 22888 11354
rect 22836 11290 22888 11296
rect 22744 11144 22796 11150
rect 22744 11086 22796 11092
rect 22848 9178 22876 11290
rect 23400 11234 23428 11494
rect 23216 11206 23428 11234
rect 23216 11098 23244 11206
rect 23492 11150 23520 11698
rect 23124 11082 23244 11098
rect 23480 11144 23532 11150
rect 23480 11086 23532 11092
rect 23112 11076 23244 11082
rect 23164 11070 23244 11076
rect 23112 11018 23164 11024
rect 22920 10908 23296 10917
rect 22976 10906 23000 10908
rect 23056 10906 23080 10908
rect 23136 10906 23160 10908
rect 23216 10906 23240 10908
rect 22976 10854 22986 10906
rect 23230 10854 23240 10906
rect 22976 10852 23000 10854
rect 23056 10852 23080 10854
rect 23136 10852 23160 10854
rect 23216 10852 23240 10854
rect 22920 10843 23296 10852
rect 22920 9820 23296 9829
rect 22976 9818 23000 9820
rect 23056 9818 23080 9820
rect 23136 9818 23160 9820
rect 23216 9818 23240 9820
rect 22976 9766 22986 9818
rect 23230 9766 23240 9818
rect 22976 9764 23000 9766
rect 23056 9764 23080 9766
rect 23136 9764 23160 9766
rect 23216 9764 23240 9766
rect 22920 9755 23296 9764
rect 23676 9722 23704 19722
rect 24860 19508 24912 19514
rect 24860 19450 24912 19456
rect 24872 18290 24900 19450
rect 25240 19174 25268 20334
rect 26160 19854 26188 20470
rect 26252 20398 26280 21830
rect 26528 20942 26556 24006
rect 26712 23594 26740 24618
rect 26804 24290 26832 25638
rect 26896 24750 26924 25774
rect 27264 24818 27292 27270
rect 27540 27130 27568 27270
rect 28920 27228 29296 27237
rect 28976 27226 29000 27228
rect 29056 27226 29080 27228
rect 29136 27226 29160 27228
rect 29216 27226 29240 27228
rect 28976 27174 28986 27226
rect 29230 27174 29240 27226
rect 28976 27172 29000 27174
rect 29056 27172 29080 27174
rect 29136 27172 29160 27174
rect 29216 27172 29240 27174
rect 28920 27163 29296 27172
rect 29380 27130 29408 27542
rect 27528 27124 27580 27130
rect 27528 27066 27580 27072
rect 29368 27124 29420 27130
rect 29368 27066 29420 27072
rect 28724 26988 28776 26994
rect 28724 26930 28776 26936
rect 27712 26920 27764 26926
rect 27712 26862 27764 26868
rect 27528 26784 27580 26790
rect 27528 26726 27580 26732
rect 27436 26444 27488 26450
rect 27436 26386 27488 26392
rect 27160 24812 27212 24818
rect 27160 24754 27212 24760
rect 27252 24812 27304 24818
rect 27252 24754 27304 24760
rect 27344 24812 27396 24818
rect 27344 24754 27396 24760
rect 26884 24744 26936 24750
rect 26884 24686 26936 24692
rect 26976 24608 27028 24614
rect 26976 24550 27028 24556
rect 26988 24410 27016 24550
rect 26976 24404 27028 24410
rect 26976 24346 27028 24352
rect 26804 24262 27108 24290
rect 26700 23588 26752 23594
rect 26700 23530 26752 23536
rect 26516 20936 26568 20942
rect 26516 20878 26568 20884
rect 26240 20392 26292 20398
rect 26240 20334 26292 20340
rect 26332 20256 26384 20262
rect 26332 20198 26384 20204
rect 26344 19854 26372 20198
rect 26148 19848 26200 19854
rect 26148 19790 26200 19796
rect 26332 19848 26384 19854
rect 26332 19790 26384 19796
rect 26160 19378 26188 19790
rect 25964 19372 26016 19378
rect 25964 19314 26016 19320
rect 26148 19372 26200 19378
rect 26148 19314 26200 19320
rect 26424 19372 26476 19378
rect 26424 19314 26476 19320
rect 25228 19168 25280 19174
rect 25228 19110 25280 19116
rect 25780 19168 25832 19174
rect 25780 19110 25832 19116
rect 24860 18284 24912 18290
rect 24860 18226 24912 18232
rect 23940 17672 23992 17678
rect 23940 17614 23992 17620
rect 23952 17202 23980 17614
rect 25044 17536 25096 17542
rect 25044 17478 25096 17484
rect 25056 17338 25084 17478
rect 25044 17332 25096 17338
rect 25044 17274 25096 17280
rect 23848 17196 23900 17202
rect 23848 17138 23900 17144
rect 23940 17196 23992 17202
rect 23940 17138 23992 17144
rect 23860 16794 23888 17138
rect 23848 16788 23900 16794
rect 23848 16730 23900 16736
rect 23848 16584 23900 16590
rect 23848 16526 23900 16532
rect 23860 16017 23888 16526
rect 23846 16008 23902 16017
rect 23846 15943 23902 15952
rect 23952 15910 23980 17138
rect 24032 16992 24084 16998
rect 24032 16934 24084 16940
rect 24044 16590 24072 16934
rect 24032 16584 24084 16590
rect 24032 16526 24084 16532
rect 23940 15904 23992 15910
rect 23940 15846 23992 15852
rect 25240 15570 25268 19110
rect 25792 18698 25820 19110
rect 25780 18692 25832 18698
rect 25780 18634 25832 18640
rect 25976 18426 26004 19314
rect 26160 18766 26188 19314
rect 26148 18760 26200 18766
rect 26148 18702 26200 18708
rect 25964 18420 26016 18426
rect 25964 18362 26016 18368
rect 26436 18086 26464 19314
rect 26424 18080 26476 18086
rect 26424 18022 26476 18028
rect 26240 17332 26292 17338
rect 26240 17274 26292 17280
rect 26252 17202 26280 17274
rect 26056 17196 26108 17202
rect 26056 17138 26108 17144
rect 26240 17196 26292 17202
rect 26240 17138 26292 17144
rect 25872 17128 25924 17134
rect 25872 17070 25924 17076
rect 25688 17060 25740 17066
rect 25688 17002 25740 17008
rect 25320 16992 25372 16998
rect 25320 16934 25372 16940
rect 25332 16522 25360 16934
rect 25700 16590 25728 17002
rect 25780 16992 25832 16998
rect 25780 16934 25832 16940
rect 25596 16584 25648 16590
rect 25596 16526 25648 16532
rect 25688 16584 25740 16590
rect 25688 16526 25740 16532
rect 25320 16516 25372 16522
rect 25320 16458 25372 16464
rect 25608 16046 25636 16526
rect 25792 16114 25820 16934
rect 25884 16794 25912 17070
rect 25872 16788 25924 16794
rect 25872 16730 25924 16736
rect 25872 16448 25924 16454
rect 25872 16390 25924 16396
rect 25884 16182 25912 16390
rect 26068 16250 26096 17138
rect 26252 17066 26280 17138
rect 26240 17060 26292 17066
rect 26240 17002 26292 17008
rect 26528 16810 26556 20878
rect 26712 20806 26740 23530
rect 26884 22568 26936 22574
rect 26884 22510 26936 22516
rect 26792 22432 26844 22438
rect 26792 22374 26844 22380
rect 26804 21486 26832 22374
rect 26792 21480 26844 21486
rect 26792 21422 26844 21428
rect 26700 20800 26752 20806
rect 26700 20742 26752 20748
rect 26608 19168 26660 19174
rect 26608 19110 26660 19116
rect 26620 18698 26648 19110
rect 26608 18692 26660 18698
rect 26608 18634 26660 18640
rect 26436 16782 26556 16810
rect 26056 16244 26108 16250
rect 26056 16186 26108 16192
rect 25872 16176 25924 16182
rect 25872 16118 25924 16124
rect 25780 16108 25832 16114
rect 25780 16050 25832 16056
rect 25596 16040 25648 16046
rect 25596 15982 25648 15988
rect 25228 15564 25280 15570
rect 25228 15506 25280 15512
rect 23940 15428 23992 15434
rect 23940 15370 23992 15376
rect 23952 15026 23980 15370
rect 23940 15020 23992 15026
rect 23940 14962 23992 14968
rect 24032 13320 24084 13326
rect 24032 13262 24084 13268
rect 24044 12986 24072 13262
rect 24032 12980 24084 12986
rect 24032 12922 24084 12928
rect 25240 12782 25268 15506
rect 25608 15502 25636 15982
rect 25596 15496 25648 15502
rect 25596 15438 25648 15444
rect 26068 15434 26096 16186
rect 26148 16108 26200 16114
rect 26148 16050 26200 16056
rect 26160 15706 26188 16050
rect 26240 15904 26292 15910
rect 26240 15846 26292 15852
rect 26148 15700 26200 15706
rect 26148 15642 26200 15648
rect 26056 15428 26108 15434
rect 26056 15370 26108 15376
rect 26252 15162 26280 15846
rect 26240 15156 26292 15162
rect 26240 15098 26292 15104
rect 26436 15026 26464 16782
rect 26516 15904 26568 15910
rect 26516 15846 26568 15852
rect 26528 15434 26556 15846
rect 26516 15428 26568 15434
rect 26516 15370 26568 15376
rect 26712 15026 26740 20742
rect 26896 17746 26924 22510
rect 26976 21344 27028 21350
rect 26976 21286 27028 21292
rect 26988 21146 27016 21286
rect 26976 21140 27028 21146
rect 26976 21082 27028 21088
rect 27080 21010 27108 24262
rect 27172 22642 27200 24754
rect 27356 22642 27384 24754
rect 27448 24290 27476 26386
rect 27540 24818 27568 26726
rect 27724 26586 27752 26862
rect 27804 26784 27856 26790
rect 27804 26726 27856 26732
rect 27816 26586 27844 26726
rect 28180 26684 28556 26693
rect 28236 26682 28260 26684
rect 28316 26682 28340 26684
rect 28396 26682 28420 26684
rect 28476 26682 28500 26684
rect 28236 26630 28246 26682
rect 28490 26630 28500 26682
rect 28236 26628 28260 26630
rect 28316 26628 28340 26630
rect 28396 26628 28420 26630
rect 28476 26628 28500 26630
rect 28180 26619 28556 26628
rect 28736 26586 28764 26930
rect 27712 26580 27764 26586
rect 27712 26522 27764 26528
rect 27804 26580 27856 26586
rect 27804 26522 27856 26528
rect 28724 26580 28776 26586
rect 28724 26522 28776 26528
rect 27724 26466 27752 26522
rect 27724 26438 27844 26466
rect 27712 26240 27764 26246
rect 27712 26182 27764 26188
rect 27724 25770 27752 26182
rect 27712 25764 27764 25770
rect 27712 25706 27764 25712
rect 27528 24812 27580 24818
rect 27528 24754 27580 24760
rect 27448 24262 27568 24290
rect 27436 23520 27488 23526
rect 27436 23462 27488 23468
rect 27160 22636 27212 22642
rect 27160 22578 27212 22584
rect 27344 22636 27396 22642
rect 27344 22578 27396 22584
rect 27068 21004 27120 21010
rect 27068 20946 27120 20952
rect 26976 20800 27028 20806
rect 26976 20742 27028 20748
rect 26988 20602 27016 20742
rect 26976 20596 27028 20602
rect 26976 20538 27028 20544
rect 26884 17740 26936 17746
rect 26884 17682 26936 17688
rect 26896 17270 26924 17682
rect 26884 17264 26936 17270
rect 26884 17206 26936 17212
rect 27080 16046 27108 20946
rect 27172 17338 27200 22578
rect 27448 22030 27476 23462
rect 27540 22098 27568 24262
rect 27620 23792 27672 23798
rect 27620 23734 27672 23740
rect 27632 23118 27660 23734
rect 27712 23656 27764 23662
rect 27712 23598 27764 23604
rect 27724 23322 27752 23598
rect 27712 23316 27764 23322
rect 27712 23258 27764 23264
rect 27620 23112 27672 23118
rect 27620 23054 27672 23060
rect 27724 22778 27752 23258
rect 27816 22930 27844 26438
rect 28920 26140 29296 26149
rect 28976 26138 29000 26140
rect 29056 26138 29080 26140
rect 29136 26138 29160 26140
rect 29216 26138 29240 26140
rect 28976 26086 28986 26138
rect 29230 26086 29240 26138
rect 28976 26084 29000 26086
rect 29056 26084 29080 26086
rect 29136 26084 29160 26086
rect 29216 26084 29240 26086
rect 28920 26075 29296 26084
rect 29380 25974 29408 27066
rect 31116 26308 31168 26314
rect 31116 26250 31168 26256
rect 31484 26308 31536 26314
rect 31484 26250 31536 26256
rect 29000 25968 29052 25974
rect 29000 25910 29052 25916
rect 29368 25968 29420 25974
rect 29368 25910 29420 25916
rect 28180 25596 28556 25605
rect 28236 25594 28260 25596
rect 28316 25594 28340 25596
rect 28396 25594 28420 25596
rect 28476 25594 28500 25596
rect 28236 25542 28246 25594
rect 28490 25542 28500 25594
rect 28236 25540 28260 25542
rect 28316 25540 28340 25542
rect 28396 25540 28420 25542
rect 28476 25540 28500 25542
rect 28180 25531 28556 25540
rect 29012 25140 29040 25910
rect 29368 25764 29420 25770
rect 29368 25706 29420 25712
rect 28828 25112 29040 25140
rect 28828 24886 28856 25112
rect 28920 25052 29296 25061
rect 28976 25050 29000 25052
rect 29056 25050 29080 25052
rect 29136 25050 29160 25052
rect 29216 25050 29240 25052
rect 28976 24998 28986 25050
rect 29230 24998 29240 25050
rect 28976 24996 29000 24998
rect 29056 24996 29080 24998
rect 29136 24996 29160 24998
rect 29216 24996 29240 24998
rect 28920 24987 29296 24996
rect 29380 24954 29408 25706
rect 29736 25220 29788 25226
rect 29736 25162 29788 25168
rect 29368 24948 29420 24954
rect 29288 24908 29368 24936
rect 28816 24880 28868 24886
rect 28816 24822 28868 24828
rect 28724 24744 28776 24750
rect 28724 24686 28776 24692
rect 28180 24508 28556 24517
rect 28236 24506 28260 24508
rect 28316 24506 28340 24508
rect 28396 24506 28420 24508
rect 28476 24506 28500 24508
rect 28236 24454 28246 24506
rect 28490 24454 28500 24506
rect 28236 24452 28260 24454
rect 28316 24452 28340 24454
rect 28396 24452 28420 24454
rect 28476 24452 28500 24454
rect 28180 24443 28556 24452
rect 28736 23730 28764 24686
rect 28828 24274 28856 24822
rect 29000 24608 29052 24614
rect 29000 24550 29052 24556
rect 29184 24608 29236 24614
rect 29184 24550 29236 24556
rect 28816 24268 28868 24274
rect 28816 24210 28868 24216
rect 29012 24138 29040 24550
rect 29196 24410 29224 24550
rect 29184 24404 29236 24410
rect 29184 24346 29236 24352
rect 29288 24274 29316 24908
rect 29368 24890 29420 24896
rect 29460 24880 29512 24886
rect 29460 24822 29512 24828
rect 29368 24812 29420 24818
rect 29368 24754 29420 24760
rect 29380 24410 29408 24754
rect 29368 24404 29420 24410
rect 29368 24346 29420 24352
rect 29276 24268 29328 24274
rect 29276 24210 29328 24216
rect 28816 24132 28868 24138
rect 28816 24074 28868 24080
rect 29000 24132 29052 24138
rect 29000 24074 29052 24080
rect 28828 23866 28856 24074
rect 28920 23964 29296 23973
rect 28976 23962 29000 23964
rect 29056 23962 29080 23964
rect 29136 23962 29160 23964
rect 29216 23962 29240 23964
rect 28976 23910 28986 23962
rect 29230 23910 29240 23962
rect 28976 23908 29000 23910
rect 29056 23908 29080 23910
rect 29136 23908 29160 23910
rect 29216 23908 29240 23910
rect 28920 23899 29296 23908
rect 28816 23860 28868 23866
rect 28816 23802 28868 23808
rect 28080 23724 28132 23730
rect 28080 23666 28132 23672
rect 28724 23724 28776 23730
rect 28724 23666 28776 23672
rect 28816 23724 28868 23730
rect 28816 23666 28868 23672
rect 29368 23724 29420 23730
rect 29368 23666 29420 23672
rect 27988 23520 28040 23526
rect 27988 23462 28040 23468
rect 28000 23050 28028 23462
rect 27988 23044 28040 23050
rect 27988 22986 28040 22992
rect 27816 22902 28028 22930
rect 27712 22772 27764 22778
rect 27712 22714 27764 22720
rect 28000 22506 28028 22902
rect 28092 22778 28120 23666
rect 28724 23520 28776 23526
rect 28724 23462 28776 23468
rect 28180 23420 28556 23429
rect 28236 23418 28260 23420
rect 28316 23418 28340 23420
rect 28396 23418 28420 23420
rect 28476 23418 28500 23420
rect 28236 23366 28246 23418
rect 28490 23366 28500 23418
rect 28236 23364 28260 23366
rect 28316 23364 28340 23366
rect 28396 23364 28420 23366
rect 28476 23364 28500 23366
rect 28180 23355 28556 23364
rect 28356 22976 28408 22982
rect 28356 22918 28408 22924
rect 28080 22772 28132 22778
rect 28080 22714 28132 22720
rect 28368 22710 28396 22918
rect 28632 22772 28684 22778
rect 28632 22714 28684 22720
rect 28356 22704 28408 22710
rect 28356 22646 28408 22652
rect 27988 22500 28040 22506
rect 27988 22442 28040 22448
rect 28180 22332 28556 22341
rect 28236 22330 28260 22332
rect 28316 22330 28340 22332
rect 28396 22330 28420 22332
rect 28476 22330 28500 22332
rect 28236 22278 28246 22330
rect 28490 22278 28500 22330
rect 28236 22276 28260 22278
rect 28316 22276 28340 22278
rect 28396 22276 28420 22278
rect 28476 22276 28500 22278
rect 28180 22267 28556 22276
rect 27528 22092 27580 22098
rect 27528 22034 27580 22040
rect 27436 22024 27488 22030
rect 27436 21966 27488 21972
rect 27436 21888 27488 21894
rect 27436 21830 27488 21836
rect 27448 21622 27476 21830
rect 27436 21616 27488 21622
rect 27436 21558 27488 21564
rect 27448 20942 27476 21558
rect 27988 21548 28040 21554
rect 27988 21490 28040 21496
rect 27436 20936 27488 20942
rect 27436 20878 27488 20884
rect 27252 20868 27304 20874
rect 27252 20810 27304 20816
rect 27896 20868 27948 20874
rect 27896 20810 27948 20816
rect 27264 20534 27292 20810
rect 27908 20602 27936 20810
rect 27896 20596 27948 20602
rect 27896 20538 27948 20544
rect 27252 20528 27304 20534
rect 27252 20470 27304 20476
rect 27264 20058 27292 20470
rect 28000 20058 28028 21490
rect 28180 21244 28556 21253
rect 28236 21242 28260 21244
rect 28316 21242 28340 21244
rect 28396 21242 28420 21244
rect 28476 21242 28500 21244
rect 28236 21190 28246 21242
rect 28490 21190 28500 21242
rect 28236 21188 28260 21190
rect 28316 21188 28340 21190
rect 28396 21188 28420 21190
rect 28476 21188 28500 21190
rect 28180 21179 28556 21188
rect 28080 21072 28132 21078
rect 28080 21014 28132 21020
rect 28092 20874 28120 21014
rect 28644 20874 28672 22714
rect 28736 22574 28764 23462
rect 28724 22568 28776 22574
rect 28724 22510 28776 22516
rect 28080 20868 28132 20874
rect 28080 20810 28132 20816
rect 28632 20868 28684 20874
rect 28632 20810 28684 20816
rect 28180 20156 28556 20165
rect 28236 20154 28260 20156
rect 28316 20154 28340 20156
rect 28396 20154 28420 20156
rect 28476 20154 28500 20156
rect 28236 20102 28246 20154
rect 28490 20102 28500 20154
rect 28236 20100 28260 20102
rect 28316 20100 28340 20102
rect 28396 20100 28420 20102
rect 28476 20100 28500 20102
rect 28180 20091 28556 20100
rect 27252 20052 27304 20058
rect 27252 19994 27304 20000
rect 27988 20052 28040 20058
rect 27988 19994 28040 20000
rect 28736 19854 28764 22510
rect 28724 19848 28776 19854
rect 28724 19790 28776 19796
rect 28828 19802 28856 23666
rect 28920 22876 29296 22885
rect 28976 22874 29000 22876
rect 29056 22874 29080 22876
rect 29136 22874 29160 22876
rect 29216 22874 29240 22876
rect 28976 22822 28986 22874
rect 29230 22822 29240 22874
rect 28976 22820 29000 22822
rect 29056 22820 29080 22822
rect 29136 22820 29160 22822
rect 29216 22820 29240 22822
rect 28920 22811 29296 22820
rect 28920 21788 29296 21797
rect 28976 21786 29000 21788
rect 29056 21786 29080 21788
rect 29136 21786 29160 21788
rect 29216 21786 29240 21788
rect 28976 21734 28986 21786
rect 29230 21734 29240 21786
rect 28976 21732 29000 21734
rect 29056 21732 29080 21734
rect 29136 21732 29160 21734
rect 29216 21732 29240 21734
rect 28920 21723 29296 21732
rect 29000 21344 29052 21350
rect 29000 21286 29052 21292
rect 29012 20942 29040 21286
rect 29000 20936 29052 20942
rect 29000 20878 29052 20884
rect 28920 20700 29296 20709
rect 28976 20698 29000 20700
rect 29056 20698 29080 20700
rect 29136 20698 29160 20700
rect 29216 20698 29240 20700
rect 28976 20646 28986 20698
rect 29230 20646 29240 20698
rect 28976 20644 29000 20646
rect 29056 20644 29080 20646
rect 29136 20644 29160 20646
rect 29216 20644 29240 20646
rect 28920 20635 29296 20644
rect 29000 20596 29052 20602
rect 29000 20538 29052 20544
rect 29012 19854 29040 20538
rect 29380 20330 29408 23666
rect 29472 21026 29500 24822
rect 29748 24750 29776 25162
rect 29736 24744 29788 24750
rect 31128 24721 31156 26250
rect 31496 25945 31524 26250
rect 31482 25936 31538 25945
rect 31482 25871 31538 25880
rect 29736 24686 29788 24692
rect 31114 24712 31170 24721
rect 29552 24064 29604 24070
rect 29552 24006 29604 24012
rect 29564 23662 29592 24006
rect 29552 23656 29604 23662
rect 29552 23598 29604 23604
rect 29748 22094 29776 24686
rect 31114 24647 31170 24656
rect 30196 24608 30248 24614
rect 30196 24550 30248 24556
rect 30840 24608 30892 24614
rect 30840 24550 30892 24556
rect 30208 23848 30236 24550
rect 30852 24070 30880 24550
rect 30840 24064 30892 24070
rect 30840 24006 30892 24012
rect 30208 23820 30328 23848
rect 30300 23730 30328 23820
rect 30288 23724 30340 23730
rect 30288 23666 30340 23672
rect 29748 22066 29868 22094
rect 29644 22024 29696 22030
rect 29644 21966 29696 21972
rect 29552 21888 29604 21894
rect 29552 21830 29604 21836
rect 29564 21690 29592 21830
rect 29552 21684 29604 21690
rect 29552 21626 29604 21632
rect 29656 21146 29684 21966
rect 29840 21486 29868 22066
rect 29828 21480 29880 21486
rect 29828 21422 29880 21428
rect 30104 21480 30156 21486
rect 30104 21422 30156 21428
rect 29644 21140 29696 21146
rect 29644 21082 29696 21088
rect 29472 21010 29592 21026
rect 29472 21004 29604 21010
rect 29472 20998 29552 21004
rect 29552 20946 29604 20952
rect 29368 20324 29420 20330
rect 29368 20266 29420 20272
rect 29380 19854 29408 20266
rect 29656 19854 29684 21082
rect 29736 21004 29788 21010
rect 29736 20946 29788 20952
rect 29000 19848 29052 19854
rect 27344 19780 27396 19786
rect 27344 19722 27396 19728
rect 27356 19378 27384 19722
rect 27988 19440 28040 19446
rect 27988 19382 28040 19388
rect 27344 19372 27396 19378
rect 27344 19314 27396 19320
rect 27528 19372 27580 19378
rect 27528 19314 27580 19320
rect 27540 18766 27568 19314
rect 28000 18970 28028 19382
rect 28736 19310 28764 19790
rect 28828 19786 28948 19802
rect 29000 19790 29052 19796
rect 29368 19848 29420 19854
rect 29368 19790 29420 19796
rect 29644 19848 29696 19854
rect 29644 19790 29696 19796
rect 28828 19780 28960 19786
rect 28828 19774 28908 19780
rect 28908 19722 28960 19728
rect 28920 19612 29296 19621
rect 28976 19610 29000 19612
rect 29056 19610 29080 19612
rect 29136 19610 29160 19612
rect 29216 19610 29240 19612
rect 28976 19558 28986 19610
rect 29230 19558 29240 19610
rect 28976 19556 29000 19558
rect 29056 19556 29080 19558
rect 29136 19556 29160 19558
rect 29216 19556 29240 19558
rect 28920 19547 29296 19556
rect 29380 19378 29408 19790
rect 29460 19712 29512 19718
rect 29460 19654 29512 19660
rect 29368 19372 29420 19378
rect 29368 19314 29420 19320
rect 28724 19304 28776 19310
rect 28724 19246 28776 19252
rect 28180 19068 28556 19077
rect 28236 19066 28260 19068
rect 28316 19066 28340 19068
rect 28396 19066 28420 19068
rect 28476 19066 28500 19068
rect 28236 19014 28246 19066
rect 28490 19014 28500 19066
rect 28236 19012 28260 19014
rect 28316 19012 28340 19014
rect 28396 19012 28420 19014
rect 28476 19012 28500 19014
rect 28180 19003 28556 19012
rect 27988 18964 28040 18970
rect 27988 18906 28040 18912
rect 27528 18760 27580 18766
rect 27528 18702 27580 18708
rect 27540 18630 27568 18702
rect 27528 18624 27580 18630
rect 27528 18566 27580 18572
rect 28000 18290 28028 18906
rect 28448 18624 28500 18630
rect 28448 18566 28500 18572
rect 28460 18426 28488 18566
rect 28448 18420 28500 18426
rect 28448 18362 28500 18368
rect 28080 18352 28132 18358
rect 28080 18294 28132 18300
rect 27988 18284 28040 18290
rect 27988 18226 28040 18232
rect 27160 17332 27212 17338
rect 27160 17274 27212 17280
rect 27620 17264 27672 17270
rect 27620 17206 27672 17212
rect 27160 16720 27212 16726
rect 27160 16662 27212 16668
rect 27172 16114 27200 16662
rect 27632 16250 27660 17206
rect 28092 17202 28120 18294
rect 28736 18290 28764 19246
rect 28920 18524 29296 18533
rect 28976 18522 29000 18524
rect 29056 18522 29080 18524
rect 29136 18522 29160 18524
rect 29216 18522 29240 18524
rect 28976 18470 28986 18522
rect 29230 18470 29240 18522
rect 28976 18468 29000 18470
rect 29056 18468 29080 18470
rect 29136 18468 29160 18470
rect 29216 18468 29240 18470
rect 28920 18459 29296 18468
rect 29380 18358 29408 19314
rect 29472 19174 29500 19654
rect 29460 19168 29512 19174
rect 29460 19110 29512 19116
rect 29368 18352 29420 18358
rect 29368 18294 29420 18300
rect 28724 18284 28776 18290
rect 28724 18226 28776 18232
rect 29748 18222 29776 20946
rect 29736 18216 29788 18222
rect 29736 18158 29788 18164
rect 29552 18148 29604 18154
rect 29552 18090 29604 18096
rect 29460 18080 29512 18086
rect 29460 18022 29512 18028
rect 28180 17980 28556 17989
rect 28236 17978 28260 17980
rect 28316 17978 28340 17980
rect 28396 17978 28420 17980
rect 28476 17978 28500 17980
rect 28236 17926 28246 17978
rect 28490 17926 28500 17978
rect 28236 17924 28260 17926
rect 28316 17924 28340 17926
rect 28396 17924 28420 17926
rect 28476 17924 28500 17926
rect 28180 17915 28556 17924
rect 29368 17740 29420 17746
rect 29368 17682 29420 17688
rect 28724 17536 28776 17542
rect 28724 17478 28776 17484
rect 28816 17536 28868 17542
rect 28816 17478 28868 17484
rect 28736 17338 28764 17478
rect 28828 17338 28856 17478
rect 28920 17436 29296 17445
rect 28976 17434 29000 17436
rect 29056 17434 29080 17436
rect 29136 17434 29160 17436
rect 29216 17434 29240 17436
rect 28976 17382 28986 17434
rect 29230 17382 29240 17434
rect 28976 17380 29000 17382
rect 29056 17380 29080 17382
rect 29136 17380 29160 17382
rect 29216 17380 29240 17382
rect 28920 17371 29296 17380
rect 29380 17338 29408 17682
rect 28724 17332 28776 17338
rect 28724 17274 28776 17280
rect 28816 17332 28868 17338
rect 28816 17274 28868 17280
rect 29184 17332 29236 17338
rect 29184 17274 29236 17280
rect 29368 17332 29420 17338
rect 29368 17274 29420 17280
rect 29092 17264 29144 17270
rect 29012 17224 29092 17252
rect 28080 17196 28132 17202
rect 28080 17138 28132 17144
rect 28180 16892 28556 16901
rect 28236 16890 28260 16892
rect 28316 16890 28340 16892
rect 28396 16890 28420 16892
rect 28476 16890 28500 16892
rect 28236 16838 28246 16890
rect 28490 16838 28500 16890
rect 28236 16836 28260 16838
rect 28316 16836 28340 16838
rect 28396 16836 28420 16838
rect 28476 16836 28500 16838
rect 28180 16827 28556 16836
rect 28632 16788 28684 16794
rect 28632 16730 28684 16736
rect 27620 16244 27672 16250
rect 27620 16186 27672 16192
rect 27160 16108 27212 16114
rect 27160 16050 27212 16056
rect 27068 16040 27120 16046
rect 27068 15982 27120 15988
rect 27896 16040 27948 16046
rect 27896 15982 27948 15988
rect 26424 15020 26476 15026
rect 26424 14962 26476 14968
rect 26700 15020 26752 15026
rect 26700 14962 26752 14968
rect 26436 14074 26464 14962
rect 26424 14068 26476 14074
rect 26424 14010 26476 14016
rect 25780 13932 25832 13938
rect 25780 13874 25832 13880
rect 26332 13932 26384 13938
rect 26332 13874 26384 13880
rect 25412 13728 25464 13734
rect 25412 13670 25464 13676
rect 25424 12986 25452 13670
rect 25792 13530 25820 13874
rect 26148 13728 26200 13734
rect 26148 13670 26200 13676
rect 25780 13524 25832 13530
rect 25780 13466 25832 13472
rect 26160 13258 26188 13670
rect 26148 13252 26200 13258
rect 26148 13194 26200 13200
rect 26344 12986 26372 13874
rect 25412 12980 25464 12986
rect 25412 12922 25464 12928
rect 26332 12980 26384 12986
rect 26332 12922 26384 12928
rect 25412 12844 25464 12850
rect 25412 12786 25464 12792
rect 23848 12776 23900 12782
rect 23848 12718 23900 12724
rect 25228 12776 25280 12782
rect 25228 12718 25280 12724
rect 23860 11898 23888 12718
rect 24676 12096 24728 12102
rect 24676 12038 24728 12044
rect 23848 11892 23900 11898
rect 23848 11834 23900 11840
rect 23860 11150 23888 11834
rect 23848 11144 23900 11150
rect 23848 11086 23900 11092
rect 24688 11014 24716 12038
rect 25240 11354 25268 12718
rect 25424 12170 25452 12786
rect 26436 12434 26464 14010
rect 26712 13938 26740 14962
rect 26700 13932 26752 13938
rect 26344 12406 26464 12434
rect 26528 13892 26700 13920
rect 25412 12164 25464 12170
rect 25412 12106 25464 12112
rect 26056 12164 26108 12170
rect 26056 12106 26108 12112
rect 25424 11801 25452 12106
rect 25410 11792 25466 11801
rect 25410 11727 25466 11736
rect 25780 11756 25832 11762
rect 25780 11698 25832 11704
rect 25596 11552 25648 11558
rect 25596 11494 25648 11500
rect 25228 11348 25280 11354
rect 25280 11308 25360 11336
rect 25228 11290 25280 11296
rect 25228 11144 25280 11150
rect 25228 11086 25280 11092
rect 24676 11008 24728 11014
rect 24676 10950 24728 10956
rect 24400 10736 24452 10742
rect 24400 10678 24452 10684
rect 23756 10260 23808 10266
rect 23756 10202 23808 10208
rect 23768 9926 23796 10202
rect 24412 10010 24440 10678
rect 24584 10124 24636 10130
rect 24584 10066 24636 10072
rect 24320 9994 24440 10010
rect 24492 10056 24544 10062
rect 24492 9998 24544 10004
rect 24308 9988 24440 9994
rect 24360 9982 24440 9988
rect 24308 9930 24360 9936
rect 23756 9920 23808 9926
rect 23756 9862 23808 9868
rect 23664 9716 23716 9722
rect 23664 9658 23716 9664
rect 23112 9580 23164 9586
rect 23112 9522 23164 9528
rect 23124 9178 23152 9522
rect 22836 9172 22888 9178
rect 22836 9114 22888 9120
rect 23112 9172 23164 9178
rect 23112 9114 23164 9120
rect 22652 9036 22704 9042
rect 22652 8978 22704 8984
rect 22744 8968 22796 8974
rect 22744 8910 22796 8916
rect 22652 8900 22704 8906
rect 22652 8842 22704 8848
rect 22100 8832 22152 8838
rect 22100 8774 22152 8780
rect 22112 8566 22140 8774
rect 22100 8560 22152 8566
rect 22100 8502 22152 8508
rect 22192 8492 22244 8498
rect 22192 8434 22244 8440
rect 22204 8378 22232 8434
rect 22112 8350 22232 8378
rect 22112 7954 22140 8350
rect 22180 8188 22556 8197
rect 22236 8186 22260 8188
rect 22316 8186 22340 8188
rect 22396 8186 22420 8188
rect 22476 8186 22500 8188
rect 22236 8134 22246 8186
rect 22490 8134 22500 8186
rect 22236 8132 22260 8134
rect 22316 8132 22340 8134
rect 22396 8132 22420 8134
rect 22476 8132 22500 8134
rect 22180 8123 22556 8132
rect 22100 7948 22152 7954
rect 22100 7890 22152 7896
rect 22112 7206 22140 7890
rect 22100 7200 22152 7206
rect 22100 7142 22152 7148
rect 22180 7100 22556 7109
rect 22236 7098 22260 7100
rect 22316 7098 22340 7100
rect 22396 7098 22420 7100
rect 22476 7098 22500 7100
rect 22236 7046 22246 7098
rect 22490 7046 22500 7098
rect 22236 7044 22260 7046
rect 22316 7044 22340 7046
rect 22396 7044 22420 7046
rect 22476 7044 22500 7046
rect 22180 7035 22556 7044
rect 22192 6928 22244 6934
rect 22192 6870 22244 6876
rect 22008 6724 22060 6730
rect 22008 6666 22060 6672
rect 22020 6390 22048 6666
rect 22008 6384 22060 6390
rect 22008 6326 22060 6332
rect 22204 6322 22232 6870
rect 22664 6458 22692 8842
rect 22756 8634 22784 8910
rect 23676 8838 23704 9658
rect 23768 8974 23796 9862
rect 24412 8974 24440 9982
rect 24504 9382 24532 9998
rect 24492 9376 24544 9382
rect 24492 9318 24544 9324
rect 24596 8974 24624 10066
rect 24688 9926 24716 10950
rect 25044 10192 25096 10198
rect 25044 10134 25096 10140
rect 24676 9920 24728 9926
rect 24676 9862 24728 9868
rect 23756 8968 23808 8974
rect 23756 8910 23808 8916
rect 24400 8968 24452 8974
rect 24400 8910 24452 8916
rect 24584 8968 24636 8974
rect 24584 8910 24636 8916
rect 22836 8832 22888 8838
rect 22836 8774 22888 8780
rect 23664 8832 23716 8838
rect 24688 8820 24716 9862
rect 25056 9674 25084 10134
rect 25056 9654 25176 9674
rect 25056 9648 25188 9654
rect 25056 9646 25136 9648
rect 25136 9590 25188 9596
rect 24952 9580 25004 9586
rect 24952 9522 25004 9528
rect 24964 9466 24992 9522
rect 25240 9466 25268 11086
rect 25332 10606 25360 11308
rect 25608 11082 25636 11494
rect 25596 11076 25648 11082
rect 25596 11018 25648 11024
rect 25792 10810 25820 11698
rect 26068 11150 26096 12106
rect 26344 11762 26372 12406
rect 26528 11830 26556 13892
rect 26700 13874 26752 13880
rect 26700 13320 26752 13326
rect 26700 13262 26752 13268
rect 26712 12918 26740 13262
rect 26700 12912 26752 12918
rect 26700 12854 26752 12860
rect 27080 12782 27108 15982
rect 27712 15904 27764 15910
rect 27712 15846 27764 15852
rect 27724 15706 27752 15846
rect 27712 15700 27764 15706
rect 27712 15642 27764 15648
rect 27528 15496 27580 15502
rect 27528 15438 27580 15444
rect 27540 15094 27568 15438
rect 27620 15360 27672 15366
rect 27620 15302 27672 15308
rect 27528 15088 27580 15094
rect 27528 15030 27580 15036
rect 27632 15026 27660 15302
rect 27908 15162 27936 15982
rect 28180 15804 28556 15813
rect 28236 15802 28260 15804
rect 28316 15802 28340 15804
rect 28396 15802 28420 15804
rect 28476 15802 28500 15804
rect 28236 15750 28246 15802
rect 28490 15750 28500 15802
rect 28236 15748 28260 15750
rect 28316 15748 28340 15750
rect 28396 15748 28420 15750
rect 28476 15748 28500 15750
rect 28180 15739 28556 15748
rect 28264 15360 28316 15366
rect 28264 15302 28316 15308
rect 27896 15156 27948 15162
rect 27896 15098 27948 15104
rect 28276 15026 28304 15302
rect 28644 15026 28672 16730
rect 28908 16584 28960 16590
rect 29012 16538 29040 17224
rect 29092 17206 29144 17212
rect 29090 16688 29146 16697
rect 29196 16658 29224 17274
rect 29472 17270 29500 18022
rect 29460 17264 29512 17270
rect 29460 17206 29512 17212
rect 29472 16794 29500 17206
rect 29460 16788 29512 16794
rect 29460 16730 29512 16736
rect 29090 16623 29092 16632
rect 29144 16623 29146 16632
rect 29184 16652 29236 16658
rect 29092 16594 29144 16600
rect 29184 16594 29236 16600
rect 28960 16532 29040 16538
rect 28908 16526 29040 16532
rect 29460 16584 29512 16590
rect 29564 16572 29592 18090
rect 29748 17746 29776 18158
rect 29736 17740 29788 17746
rect 29736 17682 29788 17688
rect 29644 17196 29696 17202
rect 29644 17138 29696 17144
rect 29512 16544 29592 16572
rect 29460 16526 29512 16532
rect 28920 16510 29040 16526
rect 28920 16348 29296 16357
rect 28976 16346 29000 16348
rect 29056 16346 29080 16348
rect 29136 16346 29160 16348
rect 29216 16346 29240 16348
rect 28976 16294 28986 16346
rect 29230 16294 29240 16346
rect 28976 16292 29000 16294
rect 29056 16292 29080 16294
rect 29136 16292 29160 16294
rect 29216 16292 29240 16294
rect 28920 16283 29296 16292
rect 28920 15260 29296 15269
rect 28976 15258 29000 15260
rect 29056 15258 29080 15260
rect 29136 15258 29160 15260
rect 29216 15258 29240 15260
rect 28976 15206 28986 15258
rect 29230 15206 29240 15258
rect 28976 15204 29000 15206
rect 29056 15204 29080 15206
rect 29136 15204 29160 15206
rect 29216 15204 29240 15206
rect 28920 15195 29296 15204
rect 27620 15020 27672 15026
rect 27620 14962 27672 14968
rect 28264 15020 28316 15026
rect 28264 14962 28316 14968
rect 28632 15020 28684 15026
rect 28632 14962 28684 14968
rect 28180 14716 28556 14725
rect 28236 14714 28260 14716
rect 28316 14714 28340 14716
rect 28396 14714 28420 14716
rect 28476 14714 28500 14716
rect 28236 14662 28246 14714
rect 28490 14662 28500 14714
rect 28236 14660 28260 14662
rect 28316 14660 28340 14662
rect 28396 14660 28420 14662
rect 28476 14660 28500 14662
rect 28180 14651 28556 14660
rect 27252 14000 27304 14006
rect 27252 13942 27304 13948
rect 27264 13530 27292 13942
rect 27344 13728 27396 13734
rect 27344 13670 27396 13676
rect 27436 13728 27488 13734
rect 27436 13670 27488 13676
rect 27896 13728 27948 13734
rect 27896 13670 27948 13676
rect 27252 13524 27304 13530
rect 27252 13466 27304 13472
rect 27356 12986 27384 13670
rect 27344 12980 27396 12986
rect 27344 12922 27396 12928
rect 27448 12850 27476 13670
rect 27908 13326 27936 13670
rect 28180 13628 28556 13637
rect 28236 13626 28260 13628
rect 28316 13626 28340 13628
rect 28396 13626 28420 13628
rect 28476 13626 28500 13628
rect 28236 13574 28246 13626
rect 28490 13574 28500 13626
rect 28236 13572 28260 13574
rect 28316 13572 28340 13574
rect 28396 13572 28420 13574
rect 28476 13572 28500 13574
rect 28180 13563 28556 13572
rect 28644 13326 28672 14962
rect 28920 14172 29296 14181
rect 28976 14170 29000 14172
rect 29056 14170 29080 14172
rect 29136 14170 29160 14172
rect 29216 14170 29240 14172
rect 28976 14118 28986 14170
rect 29230 14118 29240 14170
rect 28976 14116 29000 14118
rect 29056 14116 29080 14118
rect 29136 14116 29160 14118
rect 29216 14116 29240 14118
rect 28920 14107 29296 14116
rect 29368 13728 29420 13734
rect 29368 13670 29420 13676
rect 29380 13530 29408 13670
rect 29564 13530 29592 16544
rect 29656 13870 29684 17138
rect 29644 13864 29696 13870
rect 29644 13806 29696 13812
rect 29368 13524 29420 13530
rect 29368 13466 29420 13472
rect 29552 13524 29604 13530
rect 29552 13466 29604 13472
rect 27896 13320 27948 13326
rect 27896 13262 27948 13268
rect 28632 13320 28684 13326
rect 28632 13262 28684 13268
rect 28644 12850 28672 13262
rect 28920 13084 29296 13093
rect 28976 13082 29000 13084
rect 29056 13082 29080 13084
rect 29136 13082 29160 13084
rect 29216 13082 29240 13084
rect 28976 13030 28986 13082
rect 29230 13030 29240 13082
rect 28976 13028 29000 13030
rect 29056 13028 29080 13030
rect 29136 13028 29160 13030
rect 29216 13028 29240 13030
rect 28920 13019 29296 13028
rect 29564 12986 29592 13466
rect 29368 12980 29420 12986
rect 29368 12922 29420 12928
rect 29552 12980 29604 12986
rect 29552 12922 29604 12928
rect 27436 12844 27488 12850
rect 27436 12786 27488 12792
rect 28632 12844 28684 12850
rect 28632 12786 28684 12792
rect 27068 12776 27120 12782
rect 27068 12718 27120 12724
rect 27528 12776 27580 12782
rect 27528 12718 27580 12724
rect 27540 12306 27568 12718
rect 28180 12540 28556 12549
rect 28236 12538 28260 12540
rect 28316 12538 28340 12540
rect 28396 12538 28420 12540
rect 28476 12538 28500 12540
rect 28236 12486 28246 12538
rect 28490 12486 28500 12538
rect 28236 12484 28260 12486
rect 28316 12484 28340 12486
rect 28396 12484 28420 12486
rect 28476 12484 28500 12486
rect 28180 12475 28556 12484
rect 27528 12300 27580 12306
rect 27528 12242 27580 12248
rect 26516 11824 26568 11830
rect 26516 11766 26568 11772
rect 26332 11756 26384 11762
rect 26332 11698 26384 11704
rect 26700 11756 26752 11762
rect 26700 11698 26752 11704
rect 26424 11552 26476 11558
rect 26424 11494 26476 11500
rect 26516 11552 26568 11558
rect 26516 11494 26568 11500
rect 26056 11144 26108 11150
rect 26056 11086 26108 11092
rect 25780 10804 25832 10810
rect 25780 10746 25832 10752
rect 25320 10600 25372 10606
rect 25320 10542 25372 10548
rect 26056 10056 26108 10062
rect 26056 9998 26108 10004
rect 25688 9580 25740 9586
rect 25688 9522 25740 9528
rect 24964 9438 25268 9466
rect 24768 9376 24820 9382
rect 24768 9318 24820 9324
rect 24780 9110 24808 9318
rect 24768 9104 24820 9110
rect 24768 9046 24820 9052
rect 24860 8832 24912 8838
rect 24688 8792 24860 8820
rect 23664 8774 23716 8780
rect 24860 8774 24912 8780
rect 22744 8628 22796 8634
rect 22744 8570 22796 8576
rect 22848 8566 22876 8774
rect 22920 8732 23296 8741
rect 22976 8730 23000 8732
rect 23056 8730 23080 8732
rect 23136 8730 23160 8732
rect 23216 8730 23240 8732
rect 22976 8678 22986 8730
rect 23230 8678 23240 8730
rect 22976 8676 23000 8678
rect 23056 8676 23080 8678
rect 23136 8676 23160 8678
rect 23216 8676 23240 8678
rect 22920 8667 23296 8676
rect 22836 8560 22888 8566
rect 22836 8502 22888 8508
rect 23388 8424 23440 8430
rect 23388 8366 23440 8372
rect 22744 8356 22796 8362
rect 22744 8298 22796 8304
rect 22756 8090 22784 8298
rect 22744 8084 22796 8090
rect 22744 8026 22796 8032
rect 23400 7954 23428 8366
rect 24676 8288 24728 8294
rect 24676 8230 24728 8236
rect 22836 7948 22888 7954
rect 22836 7890 22888 7896
rect 23388 7948 23440 7954
rect 23388 7890 23440 7896
rect 22848 7342 22876 7890
rect 22920 7644 23296 7653
rect 22976 7642 23000 7644
rect 23056 7642 23080 7644
rect 23136 7642 23160 7644
rect 23216 7642 23240 7644
rect 22976 7590 22986 7642
rect 23230 7590 23240 7642
rect 22976 7588 23000 7590
rect 23056 7588 23080 7590
rect 23136 7588 23160 7590
rect 23216 7588 23240 7590
rect 22920 7579 23296 7588
rect 23400 7546 23428 7890
rect 23664 7812 23716 7818
rect 23664 7754 23716 7760
rect 23388 7540 23440 7546
rect 23388 7482 23440 7488
rect 22836 7336 22888 7342
rect 22836 7278 22888 7284
rect 22920 6556 23296 6565
rect 22976 6554 23000 6556
rect 23056 6554 23080 6556
rect 23136 6554 23160 6556
rect 23216 6554 23240 6556
rect 22976 6502 22986 6554
rect 23230 6502 23240 6554
rect 22976 6500 23000 6502
rect 23056 6500 23080 6502
rect 23136 6500 23160 6502
rect 23216 6500 23240 6502
rect 22920 6491 23296 6500
rect 22652 6452 22704 6458
rect 22652 6394 22704 6400
rect 22100 6316 22152 6322
rect 22100 6258 22152 6264
rect 22192 6316 22244 6322
rect 22192 6258 22244 6264
rect 21652 5778 21956 5794
rect 21640 5772 21968 5778
rect 21692 5766 21916 5772
rect 21640 5714 21692 5720
rect 21916 5714 21968 5720
rect 21640 5568 21692 5574
rect 21640 5510 21692 5516
rect 21652 5370 21680 5510
rect 21640 5364 21692 5370
rect 21640 5306 21692 5312
rect 22112 5234 22140 6258
rect 23676 6254 23704 7754
rect 24688 7002 24716 8230
rect 24872 7954 24900 8774
rect 24860 7948 24912 7954
rect 24860 7890 24912 7896
rect 24964 7818 24992 9438
rect 25700 9042 25728 9522
rect 26068 9382 26096 9998
rect 26056 9376 26108 9382
rect 26056 9318 26108 9324
rect 26068 9178 26096 9318
rect 26436 9178 26464 11494
rect 26528 10810 26556 11494
rect 26712 11354 26740 11698
rect 26700 11348 26752 11354
rect 26700 11290 26752 11296
rect 26792 11076 26844 11082
rect 26792 11018 26844 11024
rect 26804 10810 26832 11018
rect 26516 10804 26568 10810
rect 26516 10746 26568 10752
rect 26792 10804 26844 10810
rect 26792 10746 26844 10752
rect 27540 10606 27568 12242
rect 28920 11996 29296 12005
rect 28976 11994 29000 11996
rect 29056 11994 29080 11996
rect 29136 11994 29160 11996
rect 29216 11994 29240 11996
rect 28976 11942 28986 11994
rect 29230 11942 29240 11994
rect 28976 11940 29000 11942
rect 29056 11940 29080 11942
rect 29136 11940 29160 11942
rect 29216 11940 29240 11942
rect 28920 11931 29296 11940
rect 28080 11688 28132 11694
rect 28080 11630 28132 11636
rect 28092 11354 28120 11630
rect 28180 11452 28556 11461
rect 28236 11450 28260 11452
rect 28316 11450 28340 11452
rect 28396 11450 28420 11452
rect 28476 11450 28500 11452
rect 28236 11398 28246 11450
rect 28490 11398 28500 11450
rect 28236 11396 28260 11398
rect 28316 11396 28340 11398
rect 28396 11396 28420 11398
rect 28476 11396 28500 11398
rect 28180 11387 28556 11396
rect 28080 11348 28132 11354
rect 28080 11290 28132 11296
rect 28172 11008 28224 11014
rect 28172 10950 28224 10956
rect 28184 10810 28212 10950
rect 28920 10908 29296 10917
rect 28976 10906 29000 10908
rect 29056 10906 29080 10908
rect 29136 10906 29160 10908
rect 29216 10906 29240 10908
rect 28976 10854 28986 10906
rect 29230 10854 29240 10906
rect 28976 10852 29000 10854
rect 29056 10852 29080 10854
rect 29136 10852 29160 10854
rect 29216 10852 29240 10854
rect 28920 10843 29296 10852
rect 29380 10810 29408 12922
rect 29552 12640 29604 12646
rect 29552 12582 29604 12588
rect 29564 12442 29592 12582
rect 29552 12436 29604 12442
rect 29552 12378 29604 12384
rect 28172 10804 28224 10810
rect 28172 10746 28224 10752
rect 29368 10804 29420 10810
rect 29368 10746 29420 10752
rect 27436 10600 27488 10606
rect 27436 10542 27488 10548
rect 27528 10600 27580 10606
rect 27528 10542 27580 10548
rect 26056 9172 26108 9178
rect 26056 9114 26108 9120
rect 26424 9172 26476 9178
rect 26424 9114 26476 9120
rect 25688 9036 25740 9042
rect 25688 8978 25740 8984
rect 26608 8968 26660 8974
rect 26608 8910 26660 8916
rect 26424 8900 26476 8906
rect 26424 8842 26476 8848
rect 25780 7880 25832 7886
rect 25780 7822 25832 7828
rect 24952 7812 25004 7818
rect 24952 7754 25004 7760
rect 25792 7546 25820 7822
rect 25780 7540 25832 7546
rect 25780 7482 25832 7488
rect 25596 7404 25648 7410
rect 25596 7346 25648 7352
rect 24676 6996 24728 7002
rect 24676 6938 24728 6944
rect 24124 6792 24176 6798
rect 24124 6734 24176 6740
rect 24032 6656 24084 6662
rect 24032 6598 24084 6604
rect 23756 6452 23808 6458
rect 23756 6394 23808 6400
rect 23664 6248 23716 6254
rect 23664 6190 23716 6196
rect 23572 6112 23624 6118
rect 23572 6054 23624 6060
rect 22180 6012 22556 6021
rect 22236 6010 22260 6012
rect 22316 6010 22340 6012
rect 22396 6010 22420 6012
rect 22476 6010 22500 6012
rect 22236 5958 22246 6010
rect 22490 5958 22500 6010
rect 22236 5956 22260 5958
rect 22316 5956 22340 5958
rect 22396 5956 22420 5958
rect 22476 5956 22500 5958
rect 22180 5947 22556 5956
rect 23584 5914 23612 6054
rect 23572 5908 23624 5914
rect 23572 5850 23624 5856
rect 23676 5778 23704 6190
rect 23768 5914 23796 6394
rect 23756 5908 23808 5914
rect 23756 5850 23808 5856
rect 23664 5772 23716 5778
rect 23664 5714 23716 5720
rect 24044 5710 24072 6598
rect 24136 6458 24164 6734
rect 24688 6730 24716 6938
rect 25504 6792 25556 6798
rect 25504 6734 25556 6740
rect 24676 6724 24728 6730
rect 24676 6666 24728 6672
rect 24216 6656 24268 6662
rect 24216 6598 24268 6604
rect 24124 6452 24176 6458
rect 24124 6394 24176 6400
rect 24228 5710 24256 6598
rect 25516 6186 25544 6734
rect 25608 6390 25636 7346
rect 26436 6662 26464 8842
rect 26620 8634 26648 8910
rect 26884 8832 26936 8838
rect 26884 8774 26936 8780
rect 26608 8628 26660 8634
rect 26608 8570 26660 8576
rect 26896 8537 26924 8774
rect 27344 8628 27396 8634
rect 27344 8570 27396 8576
rect 26882 8528 26938 8537
rect 26882 8463 26938 8472
rect 27068 8424 27120 8430
rect 27068 8366 27120 8372
rect 27080 8090 27108 8366
rect 27068 8084 27120 8090
rect 27068 8026 27120 8032
rect 27356 7750 27384 8570
rect 27448 8294 27476 10542
rect 29000 10464 29052 10470
rect 29000 10406 29052 10412
rect 28180 10364 28556 10373
rect 28236 10362 28260 10364
rect 28316 10362 28340 10364
rect 28396 10362 28420 10364
rect 28476 10362 28500 10364
rect 28236 10310 28246 10362
rect 28490 10310 28500 10362
rect 28236 10308 28260 10310
rect 28316 10308 28340 10310
rect 28396 10308 28420 10310
rect 28476 10308 28500 10310
rect 28180 10299 28556 10308
rect 29012 10010 29040 10406
rect 28828 9982 29040 10010
rect 28828 9654 28856 9982
rect 29460 9920 29512 9926
rect 29460 9862 29512 9868
rect 28920 9820 29296 9829
rect 28976 9818 29000 9820
rect 29056 9818 29080 9820
rect 29136 9818 29160 9820
rect 29216 9818 29240 9820
rect 28976 9766 28986 9818
rect 29230 9766 29240 9818
rect 28976 9764 29000 9766
rect 29056 9764 29080 9766
rect 29136 9764 29160 9766
rect 29216 9764 29240 9766
rect 28920 9755 29296 9764
rect 28080 9648 28132 9654
rect 28080 9590 28132 9596
rect 28816 9648 28868 9654
rect 28816 9590 28868 9596
rect 29092 9648 29144 9654
rect 29092 9590 29144 9596
rect 28092 8362 28120 9590
rect 28816 9512 28868 9518
rect 28816 9454 28868 9460
rect 28724 9376 28776 9382
rect 28724 9318 28776 9324
rect 28180 9276 28556 9285
rect 28236 9274 28260 9276
rect 28316 9274 28340 9276
rect 28396 9274 28420 9276
rect 28476 9274 28500 9276
rect 28236 9222 28246 9274
rect 28490 9222 28500 9274
rect 28236 9220 28260 9222
rect 28316 9220 28340 9222
rect 28396 9220 28420 9222
rect 28476 9220 28500 9222
rect 28180 9211 28556 9220
rect 28736 9178 28764 9318
rect 28724 9172 28776 9178
rect 28724 9114 28776 9120
rect 28828 9042 28856 9454
rect 29104 9178 29132 9590
rect 29092 9172 29144 9178
rect 29092 9114 29144 9120
rect 28816 9036 28868 9042
rect 28816 8978 28868 8984
rect 28080 8356 28132 8362
rect 28080 8298 28132 8304
rect 27436 8288 27488 8294
rect 27436 8230 27488 8236
rect 27804 8288 27856 8294
rect 27804 8230 27856 8236
rect 27344 7744 27396 7750
rect 27344 7686 27396 7692
rect 27356 7274 27384 7686
rect 27448 7478 27476 8230
rect 27816 7546 27844 8230
rect 28180 8188 28556 8197
rect 28236 8186 28260 8188
rect 28316 8186 28340 8188
rect 28396 8186 28420 8188
rect 28476 8186 28500 8188
rect 28236 8134 28246 8186
rect 28490 8134 28500 8186
rect 28236 8132 28260 8134
rect 28316 8132 28340 8134
rect 28396 8132 28420 8134
rect 28476 8132 28500 8134
rect 28180 8123 28556 8132
rect 28828 7886 28856 8978
rect 29472 8974 29500 9862
rect 29656 9654 29684 13806
rect 29748 13190 29776 17682
rect 29840 17270 29868 21422
rect 30116 20602 30144 21422
rect 30656 21344 30708 21350
rect 30656 21286 30708 21292
rect 30668 20942 30696 21286
rect 30656 20936 30708 20942
rect 30656 20878 30708 20884
rect 31116 20868 31168 20874
rect 31116 20810 31168 20816
rect 30564 20800 30616 20806
rect 30564 20742 30616 20748
rect 31024 20800 31076 20806
rect 31024 20742 31076 20748
rect 30104 20596 30156 20602
rect 30104 20538 30156 20544
rect 30576 20466 30604 20742
rect 31036 20534 31064 20742
rect 31024 20528 31076 20534
rect 31024 20470 31076 20476
rect 30564 20460 30616 20466
rect 30564 20402 30616 20408
rect 30576 18698 30604 20402
rect 30656 19168 30708 19174
rect 30656 19110 30708 19116
rect 30564 18692 30616 18698
rect 30564 18634 30616 18640
rect 30196 17808 30248 17814
rect 30196 17750 30248 17756
rect 29920 17536 29972 17542
rect 29920 17478 29972 17484
rect 29932 17338 29960 17478
rect 29920 17332 29972 17338
rect 29920 17274 29972 17280
rect 29828 17264 29880 17270
rect 29828 17206 29880 17212
rect 29920 16788 29972 16794
rect 29920 16730 29972 16736
rect 29932 13462 29960 16730
rect 30208 16590 30236 17750
rect 30576 17202 30604 18634
rect 30564 17196 30616 17202
rect 30564 17138 30616 17144
rect 30196 16584 30248 16590
rect 30196 16526 30248 16532
rect 30668 16522 30696 19110
rect 30932 17128 30984 17134
rect 30932 17070 30984 17076
rect 30944 16697 30972 17070
rect 30930 16688 30986 16697
rect 30930 16623 30986 16632
rect 30944 16590 30972 16623
rect 30932 16584 30984 16590
rect 30932 16526 30984 16532
rect 30656 16516 30708 16522
rect 30656 16458 30708 16464
rect 30104 13864 30156 13870
rect 30104 13806 30156 13812
rect 30012 13796 30064 13802
rect 30012 13738 30064 13744
rect 29920 13456 29972 13462
rect 29920 13398 29972 13404
rect 29828 13252 29880 13258
rect 29828 13194 29880 13200
rect 29736 13184 29788 13190
rect 29736 13126 29788 13132
rect 29840 12986 29868 13194
rect 29828 12980 29880 12986
rect 29828 12922 29880 12928
rect 29736 10804 29788 10810
rect 29736 10746 29788 10752
rect 29748 10062 29776 10746
rect 29932 10266 29960 13398
rect 30024 12306 30052 13738
rect 30116 13326 30144 13806
rect 30104 13320 30156 13326
rect 30104 13262 30156 13268
rect 30668 13258 30696 16458
rect 30656 13252 30708 13258
rect 30656 13194 30708 13200
rect 30196 13184 30248 13190
rect 30196 13126 30248 13132
rect 30104 12640 30156 12646
rect 30104 12582 30156 12588
rect 30012 12300 30064 12306
rect 30012 12242 30064 12248
rect 30116 12170 30144 12582
rect 30208 12306 30236 13126
rect 30196 12300 30248 12306
rect 30196 12242 30248 12248
rect 30104 12164 30156 12170
rect 30104 12106 30156 12112
rect 30208 10826 30236 12242
rect 30116 10798 30236 10826
rect 29920 10260 29972 10266
rect 29920 10202 29972 10208
rect 30116 10130 30144 10798
rect 30196 10600 30248 10606
rect 30196 10542 30248 10548
rect 30208 10130 30236 10542
rect 30104 10124 30156 10130
rect 30104 10066 30156 10072
rect 30196 10124 30248 10130
rect 30196 10066 30248 10072
rect 29736 10056 29788 10062
rect 29736 9998 29788 10004
rect 30012 9920 30064 9926
rect 30012 9862 30064 9868
rect 30024 9722 30052 9862
rect 30208 9722 30236 10066
rect 30668 9994 30696 13194
rect 30656 9988 30708 9994
rect 30656 9930 30708 9936
rect 30748 9988 30800 9994
rect 30748 9930 30800 9936
rect 30472 9920 30524 9926
rect 30472 9862 30524 9868
rect 30484 9722 30512 9862
rect 30012 9716 30064 9722
rect 30012 9658 30064 9664
rect 30196 9716 30248 9722
rect 30196 9658 30248 9664
rect 30472 9716 30524 9722
rect 30472 9658 30524 9664
rect 29644 9648 29696 9654
rect 29644 9590 29696 9596
rect 30760 9586 30788 9930
rect 31024 9920 31076 9926
rect 31024 9862 31076 9868
rect 30748 9580 30800 9586
rect 30748 9522 30800 9528
rect 30760 9178 30788 9522
rect 30748 9172 30800 9178
rect 30748 9114 30800 9120
rect 31036 8974 31064 9862
rect 29460 8968 29512 8974
rect 29460 8910 29512 8916
rect 31024 8968 31076 8974
rect 31024 8910 31076 8916
rect 28920 8732 29296 8741
rect 28976 8730 29000 8732
rect 29056 8730 29080 8732
rect 29136 8730 29160 8732
rect 29216 8730 29240 8732
rect 28976 8678 28986 8730
rect 29230 8678 29240 8730
rect 28976 8676 29000 8678
rect 29056 8676 29080 8678
rect 29136 8676 29160 8678
rect 29216 8676 29240 8678
rect 28920 8667 29296 8676
rect 29368 8492 29420 8498
rect 29368 8434 29420 8440
rect 28816 7880 28868 7886
rect 28816 7822 28868 7828
rect 28632 7812 28684 7818
rect 28632 7754 28684 7760
rect 28644 7546 28672 7754
rect 28920 7644 29296 7653
rect 28976 7642 29000 7644
rect 29056 7642 29080 7644
rect 29136 7642 29160 7644
rect 29216 7642 29240 7644
rect 28976 7590 28986 7642
rect 29230 7590 29240 7642
rect 28976 7588 29000 7590
rect 29056 7588 29080 7590
rect 29136 7588 29160 7590
rect 29216 7588 29240 7590
rect 28920 7579 29296 7588
rect 27804 7540 27856 7546
rect 27804 7482 27856 7488
rect 28632 7540 28684 7546
rect 28632 7482 28684 7488
rect 27436 7472 27488 7478
rect 27436 7414 27488 7420
rect 27344 7268 27396 7274
rect 27344 7210 27396 7216
rect 28180 7100 28556 7109
rect 28236 7098 28260 7100
rect 28316 7098 28340 7100
rect 28396 7098 28420 7100
rect 28476 7098 28500 7100
rect 28236 7046 28246 7098
rect 28490 7046 28500 7098
rect 28236 7044 28260 7046
rect 28316 7044 28340 7046
rect 28396 7044 28420 7046
rect 28476 7044 28500 7046
rect 28180 7035 28556 7044
rect 25780 6656 25832 6662
rect 25780 6598 25832 6604
rect 26424 6656 26476 6662
rect 26424 6598 26476 6604
rect 25596 6384 25648 6390
rect 25596 6326 25648 6332
rect 25504 6180 25556 6186
rect 25504 6122 25556 6128
rect 25792 6118 25820 6598
rect 28920 6556 29296 6565
rect 28976 6554 29000 6556
rect 29056 6554 29080 6556
rect 29136 6554 29160 6556
rect 29216 6554 29240 6556
rect 28976 6502 28986 6554
rect 29230 6502 29240 6554
rect 28976 6500 29000 6502
rect 29056 6500 29080 6502
rect 29136 6500 29160 6502
rect 29216 6500 29240 6502
rect 28920 6491 29296 6500
rect 25780 6112 25832 6118
rect 25780 6054 25832 6060
rect 25792 5846 25820 6054
rect 28180 6012 28556 6021
rect 28236 6010 28260 6012
rect 28316 6010 28340 6012
rect 28396 6010 28420 6012
rect 28476 6010 28500 6012
rect 28236 5958 28246 6010
rect 28490 5958 28500 6010
rect 28236 5956 28260 5958
rect 28316 5956 28340 5958
rect 28396 5956 28420 5958
rect 28476 5956 28500 5958
rect 28180 5947 28556 5956
rect 25780 5840 25832 5846
rect 25780 5782 25832 5788
rect 24032 5704 24084 5710
rect 24032 5646 24084 5652
rect 24216 5704 24268 5710
rect 24216 5646 24268 5652
rect 22920 5468 23296 5477
rect 22976 5466 23000 5468
rect 23056 5466 23080 5468
rect 23136 5466 23160 5468
rect 23216 5466 23240 5468
rect 22976 5414 22986 5466
rect 23230 5414 23240 5466
rect 22976 5412 23000 5414
rect 23056 5412 23080 5414
rect 23136 5412 23160 5414
rect 23216 5412 23240 5414
rect 22920 5403 23296 5412
rect 28920 5468 29296 5477
rect 28976 5466 29000 5468
rect 29056 5466 29080 5468
rect 29136 5466 29160 5468
rect 29216 5466 29240 5468
rect 28976 5414 28986 5466
rect 29230 5414 29240 5466
rect 28976 5412 29000 5414
rect 29056 5412 29080 5414
rect 29136 5412 29160 5414
rect 29216 5412 29240 5414
rect 28920 5403 29296 5412
rect 22100 5228 22152 5234
rect 22100 5170 22152 5176
rect 21548 5092 21600 5098
rect 21548 5034 21600 5040
rect 21364 5024 21416 5030
rect 21364 4966 21416 4972
rect 19892 4684 19944 4690
rect 19892 4626 19944 4632
rect 21376 4622 21404 4966
rect 22112 4826 22140 5170
rect 22180 4924 22556 4933
rect 22236 4922 22260 4924
rect 22316 4922 22340 4924
rect 22396 4922 22420 4924
rect 22476 4922 22500 4924
rect 22236 4870 22246 4922
rect 22490 4870 22500 4922
rect 22236 4868 22260 4870
rect 22316 4868 22340 4870
rect 22396 4868 22420 4870
rect 22476 4868 22500 4870
rect 22180 4859 22556 4868
rect 28180 4924 28556 4933
rect 28236 4922 28260 4924
rect 28316 4922 28340 4924
rect 28396 4922 28420 4924
rect 28476 4922 28500 4924
rect 28236 4870 28246 4922
rect 28490 4870 28500 4922
rect 28236 4868 28260 4870
rect 28316 4868 28340 4870
rect 28396 4868 28420 4870
rect 28476 4868 28500 4870
rect 28180 4859 28556 4868
rect 22100 4820 22152 4826
rect 22100 4762 22152 4768
rect 18328 4616 18380 4622
rect 18328 4558 18380 4564
rect 21364 4616 21416 4622
rect 21364 4558 21416 4564
rect 16580 4548 16632 4554
rect 16580 4490 16632 4496
rect 15660 4140 15712 4146
rect 15660 4082 15712 4088
rect 15568 3936 15620 3942
rect 15568 3878 15620 3884
rect 15580 3738 15608 3878
rect 16180 3836 16556 3845
rect 16236 3834 16260 3836
rect 16316 3834 16340 3836
rect 16396 3834 16420 3836
rect 16476 3834 16500 3836
rect 16236 3782 16246 3834
rect 16490 3782 16500 3834
rect 16236 3780 16260 3782
rect 16316 3780 16340 3782
rect 16396 3780 16420 3782
rect 16476 3780 16500 3782
rect 16180 3771 16556 3780
rect 15568 3732 15620 3738
rect 15568 3674 15620 3680
rect 12164 3596 12216 3602
rect 12164 3538 12216 3544
rect 14556 3596 14608 3602
rect 14556 3538 14608 3544
rect 14648 3596 14700 3602
rect 14648 3538 14700 3544
rect 15476 3596 15528 3602
rect 15476 3538 15528 3544
rect 12440 3460 12492 3466
rect 12440 3402 12492 3408
rect 13728 3460 13780 3466
rect 13728 3402 13780 3408
rect 11888 3392 11940 3398
rect 11888 3334 11940 3340
rect 10784 3188 10836 3194
rect 10784 3130 10836 3136
rect 11612 3188 11664 3194
rect 11612 3130 11664 3136
rect 9864 3120 9916 3126
rect 9864 3062 9916 3068
rect 9772 2984 9824 2990
rect 9772 2926 9824 2932
rect 4180 2748 4556 2757
rect 4236 2746 4260 2748
rect 4316 2746 4340 2748
rect 4396 2746 4420 2748
rect 4476 2746 4500 2748
rect 4236 2694 4246 2746
rect 4490 2694 4500 2746
rect 4236 2692 4260 2694
rect 4316 2692 4340 2694
rect 4396 2692 4420 2694
rect 4476 2692 4500 2694
rect 4180 2683 4556 2692
rect 10180 2748 10556 2757
rect 10236 2746 10260 2748
rect 10316 2746 10340 2748
rect 10396 2746 10420 2748
rect 10476 2746 10500 2748
rect 10236 2694 10246 2746
rect 10490 2694 10500 2746
rect 10236 2692 10260 2694
rect 10316 2692 10340 2694
rect 10396 2692 10420 2694
rect 10476 2692 10500 2694
rect 10180 2683 10556 2692
rect 10796 2378 10824 3130
rect 11900 2446 11928 3334
rect 12452 3194 12480 3402
rect 13740 3194 13768 3402
rect 13912 3392 13964 3398
rect 13912 3334 13964 3340
rect 14096 3392 14148 3398
rect 14096 3334 14148 3340
rect 12440 3188 12492 3194
rect 12440 3130 12492 3136
rect 13728 3188 13780 3194
rect 13728 3130 13780 3136
rect 13924 2514 13952 3334
rect 14108 3194 14136 3334
rect 16592 3194 16620 4490
rect 16920 4380 17296 4389
rect 16976 4378 17000 4380
rect 17056 4378 17080 4380
rect 17136 4378 17160 4380
rect 17216 4378 17240 4380
rect 16976 4326 16986 4378
rect 17230 4326 17240 4378
rect 16976 4324 17000 4326
rect 17056 4324 17080 4326
rect 17136 4324 17160 4326
rect 17216 4324 17240 4326
rect 16920 4315 17296 4324
rect 22920 4380 23296 4389
rect 22976 4378 23000 4380
rect 23056 4378 23080 4380
rect 23136 4378 23160 4380
rect 23216 4378 23240 4380
rect 22976 4326 22986 4378
rect 23230 4326 23240 4378
rect 22976 4324 23000 4326
rect 23056 4324 23080 4326
rect 23136 4324 23160 4326
rect 23216 4324 23240 4326
rect 22920 4315 23296 4324
rect 28920 4380 29296 4389
rect 28976 4378 29000 4380
rect 29056 4378 29080 4380
rect 29136 4378 29160 4380
rect 29216 4378 29240 4380
rect 28976 4326 28986 4378
rect 29230 4326 29240 4378
rect 28976 4324 29000 4326
rect 29056 4324 29080 4326
rect 29136 4324 29160 4326
rect 29216 4324 29240 4326
rect 28920 4315 29296 4324
rect 17408 4208 17460 4214
rect 17408 4150 17460 4156
rect 17420 3738 17448 4150
rect 22180 3836 22556 3845
rect 22236 3834 22260 3836
rect 22316 3834 22340 3836
rect 22396 3834 22420 3836
rect 22476 3834 22500 3836
rect 22236 3782 22246 3834
rect 22490 3782 22500 3834
rect 22236 3780 22260 3782
rect 22316 3780 22340 3782
rect 22396 3780 22420 3782
rect 22476 3780 22500 3782
rect 22180 3771 22556 3780
rect 28180 3836 28556 3845
rect 28236 3834 28260 3836
rect 28316 3834 28340 3836
rect 28396 3834 28420 3836
rect 28476 3834 28500 3836
rect 28236 3782 28246 3834
rect 28490 3782 28500 3834
rect 28236 3780 28260 3782
rect 28316 3780 28340 3782
rect 28396 3780 28420 3782
rect 28476 3780 28500 3782
rect 28180 3771 28556 3780
rect 17408 3732 17460 3738
rect 17408 3674 17460 3680
rect 17868 3732 17920 3738
rect 17868 3674 17920 3680
rect 16672 3460 16724 3466
rect 16672 3402 16724 3408
rect 16684 3194 16712 3402
rect 16920 3292 17296 3301
rect 16976 3290 17000 3292
rect 17056 3290 17080 3292
rect 17136 3290 17160 3292
rect 17216 3290 17240 3292
rect 16976 3238 16986 3290
rect 17230 3238 17240 3290
rect 16976 3236 17000 3238
rect 17056 3236 17080 3238
rect 17136 3236 17160 3238
rect 17216 3236 17240 3238
rect 16920 3227 17296 3236
rect 14096 3188 14148 3194
rect 14096 3130 14148 3136
rect 16580 3188 16632 3194
rect 16580 3130 16632 3136
rect 16672 3188 16724 3194
rect 16672 3130 16724 3136
rect 16180 2748 16556 2757
rect 16236 2746 16260 2748
rect 16316 2746 16340 2748
rect 16396 2746 16420 2748
rect 16476 2746 16500 2748
rect 16236 2694 16246 2746
rect 16490 2694 16500 2746
rect 16236 2692 16260 2694
rect 16316 2692 16340 2694
rect 16396 2692 16420 2694
rect 16476 2692 16500 2694
rect 16180 2683 16556 2692
rect 17038 2544 17094 2553
rect 13912 2508 13964 2514
rect 17038 2479 17094 2488
rect 13912 2450 13964 2456
rect 17052 2446 17080 2479
rect 17880 2446 17908 3674
rect 22920 3292 23296 3301
rect 22976 3290 23000 3292
rect 23056 3290 23080 3292
rect 23136 3290 23160 3292
rect 23216 3290 23240 3292
rect 22976 3238 22986 3290
rect 23230 3238 23240 3290
rect 22976 3236 23000 3238
rect 23056 3236 23080 3238
rect 23136 3236 23160 3238
rect 23216 3236 23240 3238
rect 22920 3227 23296 3236
rect 28920 3292 29296 3301
rect 28976 3290 29000 3292
rect 29056 3290 29080 3292
rect 29136 3290 29160 3292
rect 29216 3290 29240 3292
rect 28976 3238 28986 3290
rect 29230 3238 29240 3290
rect 28976 3236 29000 3238
rect 29056 3236 29080 3238
rect 29136 3236 29160 3238
rect 29216 3236 29240 3238
rect 28920 3227 29296 3236
rect 22180 2748 22556 2757
rect 22236 2746 22260 2748
rect 22316 2746 22340 2748
rect 22396 2746 22420 2748
rect 22476 2746 22500 2748
rect 22236 2694 22246 2746
rect 22490 2694 22500 2746
rect 22236 2692 22260 2694
rect 22316 2692 22340 2694
rect 22396 2692 22420 2694
rect 22476 2692 22500 2694
rect 22180 2683 22556 2692
rect 28180 2748 28556 2757
rect 28236 2746 28260 2748
rect 28316 2746 28340 2748
rect 28396 2746 28420 2748
rect 28476 2746 28500 2748
rect 28236 2694 28246 2746
rect 28490 2694 28500 2746
rect 28236 2692 28260 2694
rect 28316 2692 28340 2694
rect 28396 2692 28420 2694
rect 28476 2692 28500 2694
rect 28180 2683 28556 2692
rect 29380 2650 29408 8434
rect 31128 8090 31156 20810
rect 31208 20256 31260 20262
rect 31208 20198 31260 20204
rect 31220 19854 31248 20198
rect 31852 19984 31904 19990
rect 31852 19926 31904 19932
rect 31208 19848 31260 19854
rect 31864 19825 31892 19926
rect 31208 19790 31260 19796
rect 31850 19816 31906 19825
rect 31850 19751 31906 19760
rect 31208 14816 31260 14822
rect 31208 14758 31260 14764
rect 31220 13938 31248 14758
rect 31208 13932 31260 13938
rect 31208 13874 31260 13880
rect 31484 13864 31536 13870
rect 31484 13806 31536 13812
rect 31496 13705 31524 13806
rect 31482 13696 31538 13705
rect 31482 13631 31538 13640
rect 31116 8084 31168 8090
rect 31116 8026 31168 8032
rect 31852 7812 31904 7818
rect 31852 7754 31904 7760
rect 31864 7585 31892 7754
rect 31850 7576 31906 7585
rect 31850 7511 31906 7520
rect 31208 4480 31260 4486
rect 31208 4422 31260 4428
rect 29368 2644 29420 2650
rect 29368 2586 29420 2592
rect 31220 2446 31248 4422
rect 11888 2440 11940 2446
rect 11888 2382 11940 2388
rect 17040 2440 17092 2446
rect 17040 2382 17092 2388
rect 17868 2440 17920 2446
rect 17868 2382 17920 2388
rect 29368 2440 29420 2446
rect 29368 2382 29420 2388
rect 31208 2440 31260 2446
rect 31208 2382 31260 2388
rect 20 2372 72 2378
rect 20 2314 72 2320
rect 10784 2372 10836 2378
rect 10784 2314 10836 2320
rect 32 800 60 2314
rect 5816 2304 5868 2310
rect 5816 2246 5868 2252
rect 11612 2304 11664 2310
rect 11612 2246 11664 2252
rect 17408 2304 17460 2310
rect 17408 2246 17460 2252
rect 23480 2304 23532 2310
rect 23480 2246 23532 2252
rect 4920 2204 5296 2213
rect 4976 2202 5000 2204
rect 5056 2202 5080 2204
rect 5136 2202 5160 2204
rect 5216 2202 5240 2204
rect 4976 2150 4986 2202
rect 5230 2150 5240 2202
rect 4976 2148 5000 2150
rect 5056 2148 5080 2150
rect 5136 2148 5160 2150
rect 5216 2148 5240 2150
rect 4920 2139 5296 2148
rect 5828 800 5856 2246
rect 10920 2204 11296 2213
rect 10976 2202 11000 2204
rect 11056 2202 11080 2204
rect 11136 2202 11160 2204
rect 11216 2202 11240 2204
rect 10976 2150 10986 2202
rect 11230 2150 11240 2202
rect 10976 2148 11000 2150
rect 11056 2148 11080 2150
rect 11136 2148 11160 2150
rect 11216 2148 11240 2150
rect 10920 2139 11296 2148
rect 11624 800 11652 2246
rect 16920 2204 17296 2213
rect 16976 2202 17000 2204
rect 17056 2202 17080 2204
rect 17136 2202 17160 2204
rect 17216 2202 17240 2204
rect 16976 2150 16986 2202
rect 17230 2150 17240 2202
rect 16976 2148 17000 2150
rect 17056 2148 17080 2150
rect 17136 2148 17160 2150
rect 17216 2148 17240 2150
rect 16920 2139 17296 2148
rect 17420 800 17448 2246
rect 22920 2204 23296 2213
rect 22976 2202 23000 2204
rect 23056 2202 23080 2204
rect 23136 2202 23160 2204
rect 23216 2202 23240 2204
rect 22976 2150 22986 2202
rect 23230 2150 23240 2202
rect 22976 2148 23000 2150
rect 23056 2148 23080 2150
rect 23136 2148 23160 2150
rect 23216 2148 23240 2150
rect 22920 2139 23296 2148
rect 23492 1442 23520 2246
rect 28920 2204 29296 2213
rect 28976 2202 29000 2204
rect 29056 2202 29080 2204
rect 29136 2202 29160 2204
rect 29216 2202 29240 2204
rect 28976 2150 28986 2202
rect 29230 2150 29240 2202
rect 28976 2148 29000 2150
rect 29056 2148 29080 2150
rect 29136 2148 29160 2150
rect 29216 2148 29240 2150
rect 28920 2139 29296 2148
rect 23216 1414 23520 1442
rect 23216 800 23244 1414
rect 29012 870 29132 898
rect 29012 800 29040 870
rect 18 0 74 800
rect 5814 0 5870 800
rect 11610 0 11666 800
rect 17406 0 17462 800
rect 23202 0 23258 800
rect 28998 0 29054 800
rect 29104 762 29132 870
rect 29380 762 29408 2382
rect 31392 2304 31444 2310
rect 31392 2246 31444 2252
rect 31404 1465 31432 2246
rect 31390 1456 31446 1465
rect 31390 1391 31446 1400
rect 29104 734 29408 762
<< via2 >>
rect 4920 32666 4976 32668
rect 5000 32666 5056 32668
rect 5080 32666 5136 32668
rect 5160 32666 5216 32668
rect 5240 32666 5296 32668
rect 4920 32614 4922 32666
rect 4922 32614 4974 32666
rect 4974 32614 4976 32666
rect 5000 32614 5038 32666
rect 5038 32614 5050 32666
rect 5050 32614 5056 32666
rect 5080 32614 5102 32666
rect 5102 32614 5114 32666
rect 5114 32614 5136 32666
rect 5160 32614 5166 32666
rect 5166 32614 5178 32666
rect 5178 32614 5216 32666
rect 5240 32614 5242 32666
rect 5242 32614 5294 32666
rect 5294 32614 5296 32666
rect 4920 32612 4976 32614
rect 5000 32612 5056 32614
rect 5080 32612 5136 32614
rect 5160 32612 5216 32614
rect 5240 32612 5296 32614
rect 10920 32666 10976 32668
rect 11000 32666 11056 32668
rect 11080 32666 11136 32668
rect 11160 32666 11216 32668
rect 11240 32666 11296 32668
rect 10920 32614 10922 32666
rect 10922 32614 10974 32666
rect 10974 32614 10976 32666
rect 11000 32614 11038 32666
rect 11038 32614 11050 32666
rect 11050 32614 11056 32666
rect 11080 32614 11102 32666
rect 11102 32614 11114 32666
rect 11114 32614 11136 32666
rect 11160 32614 11166 32666
rect 11166 32614 11178 32666
rect 11178 32614 11216 32666
rect 11240 32614 11242 32666
rect 11242 32614 11294 32666
rect 11294 32614 11296 32666
rect 10920 32612 10976 32614
rect 11000 32612 11056 32614
rect 11080 32612 11136 32614
rect 11160 32612 11216 32614
rect 11240 32612 11296 32614
rect 16920 32666 16976 32668
rect 17000 32666 17056 32668
rect 17080 32666 17136 32668
rect 17160 32666 17216 32668
rect 17240 32666 17296 32668
rect 16920 32614 16922 32666
rect 16922 32614 16974 32666
rect 16974 32614 16976 32666
rect 17000 32614 17038 32666
rect 17038 32614 17050 32666
rect 17050 32614 17056 32666
rect 17080 32614 17102 32666
rect 17102 32614 17114 32666
rect 17114 32614 17136 32666
rect 17160 32614 17166 32666
rect 17166 32614 17178 32666
rect 17178 32614 17216 32666
rect 17240 32614 17242 32666
rect 17242 32614 17294 32666
rect 17294 32614 17296 32666
rect 16920 32612 16976 32614
rect 17000 32612 17056 32614
rect 17080 32612 17136 32614
rect 17160 32612 17216 32614
rect 17240 32612 17296 32614
rect 22920 32666 22976 32668
rect 23000 32666 23056 32668
rect 23080 32666 23136 32668
rect 23160 32666 23216 32668
rect 23240 32666 23296 32668
rect 22920 32614 22922 32666
rect 22922 32614 22974 32666
rect 22974 32614 22976 32666
rect 23000 32614 23038 32666
rect 23038 32614 23050 32666
rect 23050 32614 23056 32666
rect 23080 32614 23102 32666
rect 23102 32614 23114 32666
rect 23114 32614 23136 32666
rect 23160 32614 23166 32666
rect 23166 32614 23178 32666
rect 23178 32614 23216 32666
rect 23240 32614 23242 32666
rect 23242 32614 23294 32666
rect 23294 32614 23296 32666
rect 22920 32612 22976 32614
rect 23000 32612 23056 32614
rect 23080 32612 23136 32614
rect 23160 32612 23216 32614
rect 23240 32612 23296 32614
rect 28920 32666 28976 32668
rect 29000 32666 29056 32668
rect 29080 32666 29136 32668
rect 29160 32666 29216 32668
rect 29240 32666 29296 32668
rect 28920 32614 28922 32666
rect 28922 32614 28974 32666
rect 28974 32614 28976 32666
rect 29000 32614 29038 32666
rect 29038 32614 29050 32666
rect 29050 32614 29056 32666
rect 29080 32614 29102 32666
rect 29102 32614 29114 32666
rect 29114 32614 29136 32666
rect 29160 32614 29166 32666
rect 29166 32614 29178 32666
rect 29178 32614 29216 32666
rect 29240 32614 29242 32666
rect 29242 32614 29294 32666
rect 29294 32614 29296 32666
rect 28920 32612 28976 32614
rect 29000 32612 29056 32614
rect 29080 32612 29136 32614
rect 29160 32612 29216 32614
rect 29240 32612 29296 32614
rect 4180 32122 4236 32124
rect 4260 32122 4316 32124
rect 4340 32122 4396 32124
rect 4420 32122 4476 32124
rect 4500 32122 4556 32124
rect 4180 32070 4182 32122
rect 4182 32070 4234 32122
rect 4234 32070 4236 32122
rect 4260 32070 4298 32122
rect 4298 32070 4310 32122
rect 4310 32070 4316 32122
rect 4340 32070 4362 32122
rect 4362 32070 4374 32122
rect 4374 32070 4396 32122
rect 4420 32070 4426 32122
rect 4426 32070 4438 32122
rect 4438 32070 4476 32122
rect 4500 32070 4502 32122
rect 4502 32070 4554 32122
rect 4554 32070 4556 32122
rect 4180 32068 4236 32070
rect 4260 32068 4316 32070
rect 4340 32068 4396 32070
rect 4420 32068 4476 32070
rect 4500 32068 4556 32070
rect 4920 31578 4976 31580
rect 5000 31578 5056 31580
rect 5080 31578 5136 31580
rect 5160 31578 5216 31580
rect 5240 31578 5296 31580
rect 4920 31526 4922 31578
rect 4922 31526 4974 31578
rect 4974 31526 4976 31578
rect 5000 31526 5038 31578
rect 5038 31526 5050 31578
rect 5050 31526 5056 31578
rect 5080 31526 5102 31578
rect 5102 31526 5114 31578
rect 5114 31526 5136 31578
rect 5160 31526 5166 31578
rect 5166 31526 5178 31578
rect 5178 31526 5216 31578
rect 5240 31526 5242 31578
rect 5242 31526 5294 31578
rect 5294 31526 5296 31578
rect 4920 31524 4976 31526
rect 5000 31524 5056 31526
rect 5080 31524 5136 31526
rect 5160 31524 5216 31526
rect 5240 31524 5296 31526
rect 4180 31034 4236 31036
rect 4260 31034 4316 31036
rect 4340 31034 4396 31036
rect 4420 31034 4476 31036
rect 4500 31034 4556 31036
rect 4180 30982 4182 31034
rect 4182 30982 4234 31034
rect 4234 30982 4236 31034
rect 4260 30982 4298 31034
rect 4298 30982 4310 31034
rect 4310 30982 4316 31034
rect 4340 30982 4362 31034
rect 4362 30982 4374 31034
rect 4374 30982 4396 31034
rect 4420 30982 4426 31034
rect 4426 30982 4438 31034
rect 4438 30982 4476 31034
rect 4500 30982 4502 31034
rect 4502 30982 4554 31034
rect 4554 30982 4556 31034
rect 4180 30980 4236 30982
rect 4260 30980 4316 30982
rect 4340 30980 4396 30982
rect 4420 30980 4476 30982
rect 4500 30980 4556 30982
rect 938 30676 940 30696
rect 940 30676 992 30696
rect 992 30676 994 30696
rect 938 30640 994 30676
rect 4920 30490 4976 30492
rect 5000 30490 5056 30492
rect 5080 30490 5136 30492
rect 5160 30490 5216 30492
rect 5240 30490 5296 30492
rect 4920 30438 4922 30490
rect 4922 30438 4974 30490
rect 4974 30438 4976 30490
rect 5000 30438 5038 30490
rect 5038 30438 5050 30490
rect 5050 30438 5056 30490
rect 5080 30438 5102 30490
rect 5102 30438 5114 30490
rect 5114 30438 5136 30490
rect 5160 30438 5166 30490
rect 5166 30438 5178 30490
rect 5178 30438 5216 30490
rect 5240 30438 5242 30490
rect 5242 30438 5294 30490
rect 5294 30438 5296 30490
rect 4920 30436 4976 30438
rect 5000 30436 5056 30438
rect 5080 30436 5136 30438
rect 5160 30436 5216 30438
rect 5240 30436 5296 30438
rect 4180 29946 4236 29948
rect 4260 29946 4316 29948
rect 4340 29946 4396 29948
rect 4420 29946 4476 29948
rect 4500 29946 4556 29948
rect 4180 29894 4182 29946
rect 4182 29894 4234 29946
rect 4234 29894 4236 29946
rect 4260 29894 4298 29946
rect 4298 29894 4310 29946
rect 4310 29894 4316 29946
rect 4340 29894 4362 29946
rect 4362 29894 4374 29946
rect 4374 29894 4396 29946
rect 4420 29894 4426 29946
rect 4426 29894 4438 29946
rect 4438 29894 4476 29946
rect 4500 29894 4502 29946
rect 4502 29894 4554 29946
rect 4554 29894 4556 29946
rect 4180 29892 4236 29894
rect 4260 29892 4316 29894
rect 4340 29892 4396 29894
rect 4420 29892 4476 29894
rect 4500 29892 4556 29894
rect 4920 29402 4976 29404
rect 5000 29402 5056 29404
rect 5080 29402 5136 29404
rect 5160 29402 5216 29404
rect 5240 29402 5296 29404
rect 4920 29350 4922 29402
rect 4922 29350 4974 29402
rect 4974 29350 4976 29402
rect 5000 29350 5038 29402
rect 5038 29350 5050 29402
rect 5050 29350 5056 29402
rect 5080 29350 5102 29402
rect 5102 29350 5114 29402
rect 5114 29350 5136 29402
rect 5160 29350 5166 29402
rect 5166 29350 5178 29402
rect 5178 29350 5216 29402
rect 5240 29350 5242 29402
rect 5242 29350 5294 29402
rect 5294 29350 5296 29402
rect 4920 29348 4976 29350
rect 5000 29348 5056 29350
rect 5080 29348 5136 29350
rect 5160 29348 5216 29350
rect 5240 29348 5296 29350
rect 4180 28858 4236 28860
rect 4260 28858 4316 28860
rect 4340 28858 4396 28860
rect 4420 28858 4476 28860
rect 4500 28858 4556 28860
rect 4180 28806 4182 28858
rect 4182 28806 4234 28858
rect 4234 28806 4236 28858
rect 4260 28806 4298 28858
rect 4298 28806 4310 28858
rect 4310 28806 4316 28858
rect 4340 28806 4362 28858
rect 4362 28806 4374 28858
rect 4374 28806 4396 28858
rect 4420 28806 4426 28858
rect 4426 28806 4438 28858
rect 4438 28806 4476 28858
rect 4500 28806 4502 28858
rect 4502 28806 4554 28858
rect 4554 28806 4556 28858
rect 4180 28804 4236 28806
rect 4260 28804 4316 28806
rect 4340 28804 4396 28806
rect 4420 28804 4476 28806
rect 4500 28804 4556 28806
rect 4920 28314 4976 28316
rect 5000 28314 5056 28316
rect 5080 28314 5136 28316
rect 5160 28314 5216 28316
rect 5240 28314 5296 28316
rect 4920 28262 4922 28314
rect 4922 28262 4974 28314
rect 4974 28262 4976 28314
rect 5000 28262 5038 28314
rect 5038 28262 5050 28314
rect 5050 28262 5056 28314
rect 5080 28262 5102 28314
rect 5102 28262 5114 28314
rect 5114 28262 5136 28314
rect 5160 28262 5166 28314
rect 5166 28262 5178 28314
rect 5178 28262 5216 28314
rect 5240 28262 5242 28314
rect 5242 28262 5294 28314
rect 5294 28262 5296 28314
rect 4920 28260 4976 28262
rect 5000 28260 5056 28262
rect 5080 28260 5136 28262
rect 5160 28260 5216 28262
rect 5240 28260 5296 28262
rect 4180 27770 4236 27772
rect 4260 27770 4316 27772
rect 4340 27770 4396 27772
rect 4420 27770 4476 27772
rect 4500 27770 4556 27772
rect 4180 27718 4182 27770
rect 4182 27718 4234 27770
rect 4234 27718 4236 27770
rect 4260 27718 4298 27770
rect 4298 27718 4310 27770
rect 4310 27718 4316 27770
rect 4340 27718 4362 27770
rect 4362 27718 4374 27770
rect 4374 27718 4396 27770
rect 4420 27718 4426 27770
rect 4426 27718 4438 27770
rect 4438 27718 4476 27770
rect 4500 27718 4502 27770
rect 4502 27718 4554 27770
rect 4554 27718 4556 27770
rect 4180 27716 4236 27718
rect 4260 27716 4316 27718
rect 4340 27716 4396 27718
rect 4420 27716 4476 27718
rect 4500 27716 4556 27718
rect 4180 26682 4236 26684
rect 4260 26682 4316 26684
rect 4340 26682 4396 26684
rect 4420 26682 4476 26684
rect 4500 26682 4556 26684
rect 4180 26630 4182 26682
rect 4182 26630 4234 26682
rect 4234 26630 4236 26682
rect 4260 26630 4298 26682
rect 4298 26630 4310 26682
rect 4310 26630 4316 26682
rect 4340 26630 4362 26682
rect 4362 26630 4374 26682
rect 4374 26630 4396 26682
rect 4420 26630 4426 26682
rect 4426 26630 4438 26682
rect 4438 26630 4476 26682
rect 4500 26630 4502 26682
rect 4502 26630 4554 26682
rect 4554 26630 4556 26682
rect 4180 26628 4236 26630
rect 4260 26628 4316 26630
rect 4340 26628 4396 26630
rect 4420 26628 4476 26630
rect 4500 26628 4556 26630
rect 938 24520 994 24576
rect 938 18400 994 18456
rect 4920 27226 4976 27228
rect 5000 27226 5056 27228
rect 5080 27226 5136 27228
rect 5160 27226 5216 27228
rect 5240 27226 5296 27228
rect 4920 27174 4922 27226
rect 4922 27174 4974 27226
rect 4974 27174 4976 27226
rect 5000 27174 5038 27226
rect 5038 27174 5050 27226
rect 5050 27174 5056 27226
rect 5080 27174 5102 27226
rect 5102 27174 5114 27226
rect 5114 27174 5136 27226
rect 5160 27174 5166 27226
rect 5166 27174 5178 27226
rect 5178 27174 5216 27226
rect 5240 27174 5242 27226
rect 5242 27174 5294 27226
rect 5294 27174 5296 27226
rect 4920 27172 4976 27174
rect 5000 27172 5056 27174
rect 5080 27172 5136 27174
rect 5160 27172 5216 27174
rect 5240 27172 5296 27174
rect 4920 26138 4976 26140
rect 5000 26138 5056 26140
rect 5080 26138 5136 26140
rect 5160 26138 5216 26140
rect 5240 26138 5296 26140
rect 4920 26086 4922 26138
rect 4922 26086 4974 26138
rect 4974 26086 4976 26138
rect 5000 26086 5038 26138
rect 5038 26086 5050 26138
rect 5050 26086 5056 26138
rect 5080 26086 5102 26138
rect 5102 26086 5114 26138
rect 5114 26086 5136 26138
rect 5160 26086 5166 26138
rect 5166 26086 5178 26138
rect 5178 26086 5216 26138
rect 5240 26086 5242 26138
rect 5242 26086 5294 26138
rect 5294 26086 5296 26138
rect 4920 26084 4976 26086
rect 5000 26084 5056 26086
rect 5080 26084 5136 26086
rect 5160 26084 5216 26086
rect 5240 26084 5296 26086
rect 4180 25594 4236 25596
rect 4260 25594 4316 25596
rect 4340 25594 4396 25596
rect 4420 25594 4476 25596
rect 4500 25594 4556 25596
rect 4180 25542 4182 25594
rect 4182 25542 4234 25594
rect 4234 25542 4236 25594
rect 4260 25542 4298 25594
rect 4298 25542 4310 25594
rect 4310 25542 4316 25594
rect 4340 25542 4362 25594
rect 4362 25542 4374 25594
rect 4374 25542 4396 25594
rect 4420 25542 4426 25594
rect 4426 25542 4438 25594
rect 4438 25542 4476 25594
rect 4500 25542 4502 25594
rect 4502 25542 4554 25594
rect 4554 25542 4556 25594
rect 4180 25540 4236 25542
rect 4260 25540 4316 25542
rect 4340 25540 4396 25542
rect 4420 25540 4476 25542
rect 4500 25540 4556 25542
rect 4180 24506 4236 24508
rect 4260 24506 4316 24508
rect 4340 24506 4396 24508
rect 4420 24506 4476 24508
rect 4500 24506 4556 24508
rect 4180 24454 4182 24506
rect 4182 24454 4234 24506
rect 4234 24454 4236 24506
rect 4260 24454 4298 24506
rect 4298 24454 4310 24506
rect 4310 24454 4316 24506
rect 4340 24454 4362 24506
rect 4362 24454 4374 24506
rect 4374 24454 4396 24506
rect 4420 24454 4426 24506
rect 4426 24454 4438 24506
rect 4438 24454 4476 24506
rect 4500 24454 4502 24506
rect 4502 24454 4554 24506
rect 4554 24454 4556 24506
rect 4180 24452 4236 24454
rect 4260 24452 4316 24454
rect 4340 24452 4396 24454
rect 4420 24452 4476 24454
rect 4500 24452 4556 24454
rect 4180 23418 4236 23420
rect 4260 23418 4316 23420
rect 4340 23418 4396 23420
rect 4420 23418 4476 23420
rect 4500 23418 4556 23420
rect 4180 23366 4182 23418
rect 4182 23366 4234 23418
rect 4234 23366 4236 23418
rect 4260 23366 4298 23418
rect 4298 23366 4310 23418
rect 4310 23366 4316 23418
rect 4340 23366 4362 23418
rect 4362 23366 4374 23418
rect 4374 23366 4396 23418
rect 4420 23366 4426 23418
rect 4426 23366 4438 23418
rect 4438 23366 4476 23418
rect 4500 23366 4502 23418
rect 4502 23366 4554 23418
rect 4554 23366 4556 23418
rect 4180 23364 4236 23366
rect 4260 23364 4316 23366
rect 4340 23364 4396 23366
rect 4420 23364 4476 23366
rect 4500 23364 4556 23366
rect 4920 25050 4976 25052
rect 5000 25050 5056 25052
rect 5080 25050 5136 25052
rect 5160 25050 5216 25052
rect 5240 25050 5296 25052
rect 4920 24998 4922 25050
rect 4922 24998 4974 25050
rect 4974 24998 4976 25050
rect 5000 24998 5038 25050
rect 5038 24998 5050 25050
rect 5050 24998 5056 25050
rect 5080 24998 5102 25050
rect 5102 24998 5114 25050
rect 5114 24998 5136 25050
rect 5160 24998 5166 25050
rect 5166 24998 5178 25050
rect 5178 24998 5216 25050
rect 5240 24998 5242 25050
rect 5242 24998 5294 25050
rect 5294 24998 5296 25050
rect 4920 24996 4976 24998
rect 5000 24996 5056 24998
rect 5080 24996 5136 24998
rect 5160 24996 5216 24998
rect 5240 24996 5296 24998
rect 4920 23962 4976 23964
rect 5000 23962 5056 23964
rect 5080 23962 5136 23964
rect 5160 23962 5216 23964
rect 5240 23962 5296 23964
rect 4920 23910 4922 23962
rect 4922 23910 4974 23962
rect 4974 23910 4976 23962
rect 5000 23910 5038 23962
rect 5038 23910 5050 23962
rect 5050 23910 5056 23962
rect 5080 23910 5102 23962
rect 5102 23910 5114 23962
rect 5114 23910 5136 23962
rect 5160 23910 5166 23962
rect 5166 23910 5178 23962
rect 5178 23910 5216 23962
rect 5240 23910 5242 23962
rect 5242 23910 5294 23962
rect 5294 23910 5296 23962
rect 4920 23908 4976 23910
rect 5000 23908 5056 23910
rect 5080 23908 5136 23910
rect 5160 23908 5216 23910
rect 5240 23908 5296 23910
rect 4180 22330 4236 22332
rect 4260 22330 4316 22332
rect 4340 22330 4396 22332
rect 4420 22330 4476 22332
rect 4500 22330 4556 22332
rect 4180 22278 4182 22330
rect 4182 22278 4234 22330
rect 4234 22278 4236 22330
rect 4260 22278 4298 22330
rect 4298 22278 4310 22330
rect 4310 22278 4316 22330
rect 4340 22278 4362 22330
rect 4362 22278 4374 22330
rect 4374 22278 4396 22330
rect 4420 22278 4426 22330
rect 4426 22278 4438 22330
rect 4438 22278 4476 22330
rect 4500 22278 4502 22330
rect 4502 22278 4554 22330
rect 4554 22278 4556 22330
rect 4180 22276 4236 22278
rect 4260 22276 4316 22278
rect 4340 22276 4396 22278
rect 4420 22276 4476 22278
rect 4500 22276 4556 22278
rect 4180 21242 4236 21244
rect 4260 21242 4316 21244
rect 4340 21242 4396 21244
rect 4420 21242 4476 21244
rect 4500 21242 4556 21244
rect 4180 21190 4182 21242
rect 4182 21190 4234 21242
rect 4234 21190 4236 21242
rect 4260 21190 4298 21242
rect 4298 21190 4310 21242
rect 4310 21190 4316 21242
rect 4340 21190 4362 21242
rect 4362 21190 4374 21242
rect 4374 21190 4396 21242
rect 4420 21190 4426 21242
rect 4426 21190 4438 21242
rect 4438 21190 4476 21242
rect 4500 21190 4502 21242
rect 4502 21190 4554 21242
rect 4554 21190 4556 21242
rect 4180 21188 4236 21190
rect 4260 21188 4316 21190
rect 4340 21188 4396 21190
rect 4420 21188 4476 21190
rect 4500 21188 4556 21190
rect 4180 20154 4236 20156
rect 4260 20154 4316 20156
rect 4340 20154 4396 20156
rect 4420 20154 4476 20156
rect 4500 20154 4556 20156
rect 4180 20102 4182 20154
rect 4182 20102 4234 20154
rect 4234 20102 4236 20154
rect 4260 20102 4298 20154
rect 4298 20102 4310 20154
rect 4310 20102 4316 20154
rect 4340 20102 4362 20154
rect 4362 20102 4374 20154
rect 4374 20102 4396 20154
rect 4420 20102 4426 20154
rect 4426 20102 4438 20154
rect 4438 20102 4476 20154
rect 4500 20102 4502 20154
rect 4502 20102 4554 20154
rect 4554 20102 4556 20154
rect 4180 20100 4236 20102
rect 4260 20100 4316 20102
rect 4340 20100 4396 20102
rect 4420 20100 4476 20102
rect 4500 20100 4556 20102
rect 1490 12280 1546 12336
rect 4180 19066 4236 19068
rect 4260 19066 4316 19068
rect 4340 19066 4396 19068
rect 4420 19066 4476 19068
rect 4500 19066 4556 19068
rect 4180 19014 4182 19066
rect 4182 19014 4234 19066
rect 4234 19014 4236 19066
rect 4260 19014 4298 19066
rect 4298 19014 4310 19066
rect 4310 19014 4316 19066
rect 4340 19014 4362 19066
rect 4362 19014 4374 19066
rect 4374 19014 4396 19066
rect 4420 19014 4426 19066
rect 4426 19014 4438 19066
rect 4438 19014 4476 19066
rect 4500 19014 4502 19066
rect 4502 19014 4554 19066
rect 4554 19014 4556 19066
rect 4180 19012 4236 19014
rect 4260 19012 4316 19014
rect 4340 19012 4396 19014
rect 4420 19012 4476 19014
rect 4500 19012 4556 19014
rect 4920 22874 4976 22876
rect 5000 22874 5056 22876
rect 5080 22874 5136 22876
rect 5160 22874 5216 22876
rect 5240 22874 5296 22876
rect 4920 22822 4922 22874
rect 4922 22822 4974 22874
rect 4974 22822 4976 22874
rect 5000 22822 5038 22874
rect 5038 22822 5050 22874
rect 5050 22822 5056 22874
rect 5080 22822 5102 22874
rect 5102 22822 5114 22874
rect 5114 22822 5136 22874
rect 5160 22822 5166 22874
rect 5166 22822 5178 22874
rect 5178 22822 5216 22874
rect 5240 22822 5242 22874
rect 5242 22822 5294 22874
rect 5294 22822 5296 22874
rect 4920 22820 4976 22822
rect 5000 22820 5056 22822
rect 5080 22820 5136 22822
rect 5160 22820 5216 22822
rect 5240 22820 5296 22822
rect 4920 21786 4976 21788
rect 5000 21786 5056 21788
rect 5080 21786 5136 21788
rect 5160 21786 5216 21788
rect 5240 21786 5296 21788
rect 4920 21734 4922 21786
rect 4922 21734 4974 21786
rect 4974 21734 4976 21786
rect 5000 21734 5038 21786
rect 5038 21734 5050 21786
rect 5050 21734 5056 21786
rect 5080 21734 5102 21786
rect 5102 21734 5114 21786
rect 5114 21734 5136 21786
rect 5160 21734 5166 21786
rect 5166 21734 5178 21786
rect 5178 21734 5216 21786
rect 5240 21734 5242 21786
rect 5242 21734 5294 21786
rect 5294 21734 5296 21786
rect 4920 21732 4976 21734
rect 5000 21732 5056 21734
rect 5080 21732 5136 21734
rect 5160 21732 5216 21734
rect 5240 21732 5296 21734
rect 4920 20698 4976 20700
rect 5000 20698 5056 20700
rect 5080 20698 5136 20700
rect 5160 20698 5216 20700
rect 5240 20698 5296 20700
rect 4920 20646 4922 20698
rect 4922 20646 4974 20698
rect 4974 20646 4976 20698
rect 5000 20646 5038 20698
rect 5038 20646 5050 20698
rect 5050 20646 5056 20698
rect 5080 20646 5102 20698
rect 5102 20646 5114 20698
rect 5114 20646 5136 20698
rect 5160 20646 5166 20698
rect 5166 20646 5178 20698
rect 5178 20646 5216 20698
rect 5240 20646 5242 20698
rect 5242 20646 5294 20698
rect 5294 20646 5296 20698
rect 4920 20644 4976 20646
rect 5000 20644 5056 20646
rect 5080 20644 5136 20646
rect 5160 20644 5216 20646
rect 5240 20644 5296 20646
rect 4180 17978 4236 17980
rect 4260 17978 4316 17980
rect 4340 17978 4396 17980
rect 4420 17978 4476 17980
rect 4500 17978 4556 17980
rect 4180 17926 4182 17978
rect 4182 17926 4234 17978
rect 4234 17926 4236 17978
rect 4260 17926 4298 17978
rect 4298 17926 4310 17978
rect 4310 17926 4316 17978
rect 4340 17926 4362 17978
rect 4362 17926 4374 17978
rect 4374 17926 4396 17978
rect 4420 17926 4426 17978
rect 4426 17926 4438 17978
rect 4438 17926 4476 17978
rect 4500 17926 4502 17978
rect 4502 17926 4554 17978
rect 4554 17926 4556 17978
rect 4180 17924 4236 17926
rect 4260 17924 4316 17926
rect 4340 17924 4396 17926
rect 4420 17924 4476 17926
rect 4500 17924 4556 17926
rect 4180 16890 4236 16892
rect 4260 16890 4316 16892
rect 4340 16890 4396 16892
rect 4420 16890 4476 16892
rect 4500 16890 4556 16892
rect 4180 16838 4182 16890
rect 4182 16838 4234 16890
rect 4234 16838 4236 16890
rect 4260 16838 4298 16890
rect 4298 16838 4310 16890
rect 4310 16838 4316 16890
rect 4340 16838 4362 16890
rect 4362 16838 4374 16890
rect 4374 16838 4396 16890
rect 4420 16838 4426 16890
rect 4426 16838 4438 16890
rect 4438 16838 4476 16890
rect 4500 16838 4502 16890
rect 4502 16838 4554 16890
rect 4554 16838 4556 16890
rect 4180 16836 4236 16838
rect 4260 16836 4316 16838
rect 4340 16836 4396 16838
rect 4420 16836 4476 16838
rect 4500 16836 4556 16838
rect 4920 19610 4976 19612
rect 5000 19610 5056 19612
rect 5080 19610 5136 19612
rect 5160 19610 5216 19612
rect 5240 19610 5296 19612
rect 4920 19558 4922 19610
rect 4922 19558 4974 19610
rect 4974 19558 4976 19610
rect 5000 19558 5038 19610
rect 5038 19558 5050 19610
rect 5050 19558 5056 19610
rect 5080 19558 5102 19610
rect 5102 19558 5114 19610
rect 5114 19558 5136 19610
rect 5160 19558 5166 19610
rect 5166 19558 5178 19610
rect 5178 19558 5216 19610
rect 5240 19558 5242 19610
rect 5242 19558 5294 19610
rect 5294 19558 5296 19610
rect 4920 19556 4976 19558
rect 5000 19556 5056 19558
rect 5080 19556 5136 19558
rect 5160 19556 5216 19558
rect 5240 19556 5296 19558
rect 10180 32122 10236 32124
rect 10260 32122 10316 32124
rect 10340 32122 10396 32124
rect 10420 32122 10476 32124
rect 10500 32122 10556 32124
rect 10180 32070 10182 32122
rect 10182 32070 10234 32122
rect 10234 32070 10236 32122
rect 10260 32070 10298 32122
rect 10298 32070 10310 32122
rect 10310 32070 10316 32122
rect 10340 32070 10362 32122
rect 10362 32070 10374 32122
rect 10374 32070 10396 32122
rect 10420 32070 10426 32122
rect 10426 32070 10438 32122
rect 10438 32070 10476 32122
rect 10500 32070 10502 32122
rect 10502 32070 10554 32122
rect 10554 32070 10556 32122
rect 10180 32068 10236 32070
rect 10260 32068 10316 32070
rect 10340 32068 10396 32070
rect 10420 32068 10476 32070
rect 10500 32068 10556 32070
rect 10920 31578 10976 31580
rect 11000 31578 11056 31580
rect 11080 31578 11136 31580
rect 11160 31578 11216 31580
rect 11240 31578 11296 31580
rect 10920 31526 10922 31578
rect 10922 31526 10974 31578
rect 10974 31526 10976 31578
rect 11000 31526 11038 31578
rect 11038 31526 11050 31578
rect 11050 31526 11056 31578
rect 11080 31526 11102 31578
rect 11102 31526 11114 31578
rect 11114 31526 11136 31578
rect 11160 31526 11166 31578
rect 11166 31526 11178 31578
rect 11178 31526 11216 31578
rect 11240 31526 11242 31578
rect 11242 31526 11294 31578
rect 11294 31526 11296 31578
rect 10920 31524 10976 31526
rect 11000 31524 11056 31526
rect 11080 31524 11136 31526
rect 11160 31524 11216 31526
rect 11240 31524 11296 31526
rect 10180 31034 10236 31036
rect 10260 31034 10316 31036
rect 10340 31034 10396 31036
rect 10420 31034 10476 31036
rect 10500 31034 10556 31036
rect 10180 30982 10182 31034
rect 10182 30982 10234 31034
rect 10234 30982 10236 31034
rect 10260 30982 10298 31034
rect 10298 30982 10310 31034
rect 10310 30982 10316 31034
rect 10340 30982 10362 31034
rect 10362 30982 10374 31034
rect 10374 30982 10396 31034
rect 10420 30982 10426 31034
rect 10426 30982 10438 31034
rect 10438 30982 10476 31034
rect 10500 30982 10502 31034
rect 10502 30982 10554 31034
rect 10554 30982 10556 31034
rect 10180 30980 10236 30982
rect 10260 30980 10316 30982
rect 10340 30980 10396 30982
rect 10420 30980 10476 30982
rect 10500 30980 10556 30982
rect 16180 32122 16236 32124
rect 16260 32122 16316 32124
rect 16340 32122 16396 32124
rect 16420 32122 16476 32124
rect 16500 32122 16556 32124
rect 16180 32070 16182 32122
rect 16182 32070 16234 32122
rect 16234 32070 16236 32122
rect 16260 32070 16298 32122
rect 16298 32070 16310 32122
rect 16310 32070 16316 32122
rect 16340 32070 16362 32122
rect 16362 32070 16374 32122
rect 16374 32070 16396 32122
rect 16420 32070 16426 32122
rect 16426 32070 16438 32122
rect 16438 32070 16476 32122
rect 16500 32070 16502 32122
rect 16502 32070 16554 32122
rect 16554 32070 16556 32122
rect 16180 32068 16236 32070
rect 16260 32068 16316 32070
rect 16340 32068 16396 32070
rect 16420 32068 16476 32070
rect 16500 32068 16556 32070
rect 10180 29946 10236 29948
rect 10260 29946 10316 29948
rect 10340 29946 10396 29948
rect 10420 29946 10476 29948
rect 10500 29946 10556 29948
rect 10180 29894 10182 29946
rect 10182 29894 10234 29946
rect 10234 29894 10236 29946
rect 10260 29894 10298 29946
rect 10298 29894 10310 29946
rect 10310 29894 10316 29946
rect 10340 29894 10362 29946
rect 10362 29894 10374 29946
rect 10374 29894 10396 29946
rect 10420 29894 10426 29946
rect 10426 29894 10438 29946
rect 10438 29894 10476 29946
rect 10500 29894 10502 29946
rect 10502 29894 10554 29946
rect 10554 29894 10556 29946
rect 10180 29892 10236 29894
rect 10260 29892 10316 29894
rect 10340 29892 10396 29894
rect 10420 29892 10476 29894
rect 10500 29892 10556 29894
rect 10180 28858 10236 28860
rect 10260 28858 10316 28860
rect 10340 28858 10396 28860
rect 10420 28858 10476 28860
rect 10500 28858 10556 28860
rect 10180 28806 10182 28858
rect 10182 28806 10234 28858
rect 10234 28806 10236 28858
rect 10260 28806 10298 28858
rect 10298 28806 10310 28858
rect 10310 28806 10316 28858
rect 10340 28806 10362 28858
rect 10362 28806 10374 28858
rect 10374 28806 10396 28858
rect 10420 28806 10426 28858
rect 10426 28806 10438 28858
rect 10438 28806 10476 28858
rect 10500 28806 10502 28858
rect 10502 28806 10554 28858
rect 10554 28806 10556 28858
rect 10180 28804 10236 28806
rect 10260 28804 10316 28806
rect 10340 28804 10396 28806
rect 10420 28804 10476 28806
rect 10500 28804 10556 28806
rect 4920 18522 4976 18524
rect 5000 18522 5056 18524
rect 5080 18522 5136 18524
rect 5160 18522 5216 18524
rect 5240 18522 5296 18524
rect 4920 18470 4922 18522
rect 4922 18470 4974 18522
rect 4974 18470 4976 18522
rect 5000 18470 5038 18522
rect 5038 18470 5050 18522
rect 5050 18470 5056 18522
rect 5080 18470 5102 18522
rect 5102 18470 5114 18522
rect 5114 18470 5136 18522
rect 5160 18470 5166 18522
rect 5166 18470 5178 18522
rect 5178 18470 5216 18522
rect 5240 18470 5242 18522
rect 5242 18470 5294 18522
rect 5294 18470 5296 18522
rect 4920 18468 4976 18470
rect 5000 18468 5056 18470
rect 5080 18468 5136 18470
rect 5160 18468 5216 18470
rect 5240 18468 5296 18470
rect 4920 17434 4976 17436
rect 5000 17434 5056 17436
rect 5080 17434 5136 17436
rect 5160 17434 5216 17436
rect 5240 17434 5296 17436
rect 4920 17382 4922 17434
rect 4922 17382 4974 17434
rect 4974 17382 4976 17434
rect 5000 17382 5038 17434
rect 5038 17382 5050 17434
rect 5050 17382 5056 17434
rect 5080 17382 5102 17434
rect 5102 17382 5114 17434
rect 5114 17382 5136 17434
rect 5160 17382 5166 17434
rect 5166 17382 5178 17434
rect 5178 17382 5216 17434
rect 5240 17382 5242 17434
rect 5242 17382 5294 17434
rect 5294 17382 5296 17434
rect 4920 17380 4976 17382
rect 5000 17380 5056 17382
rect 5080 17380 5136 17382
rect 5160 17380 5216 17382
rect 5240 17380 5296 17382
rect 4180 15802 4236 15804
rect 4260 15802 4316 15804
rect 4340 15802 4396 15804
rect 4420 15802 4476 15804
rect 4500 15802 4556 15804
rect 4180 15750 4182 15802
rect 4182 15750 4234 15802
rect 4234 15750 4236 15802
rect 4260 15750 4298 15802
rect 4298 15750 4310 15802
rect 4310 15750 4316 15802
rect 4340 15750 4362 15802
rect 4362 15750 4374 15802
rect 4374 15750 4396 15802
rect 4420 15750 4426 15802
rect 4426 15750 4438 15802
rect 4438 15750 4476 15802
rect 4500 15750 4502 15802
rect 4502 15750 4554 15802
rect 4554 15750 4556 15802
rect 4180 15748 4236 15750
rect 4260 15748 4316 15750
rect 4340 15748 4396 15750
rect 4420 15748 4476 15750
rect 4500 15748 4556 15750
rect 4180 14714 4236 14716
rect 4260 14714 4316 14716
rect 4340 14714 4396 14716
rect 4420 14714 4476 14716
rect 4500 14714 4556 14716
rect 4180 14662 4182 14714
rect 4182 14662 4234 14714
rect 4234 14662 4236 14714
rect 4260 14662 4298 14714
rect 4298 14662 4310 14714
rect 4310 14662 4316 14714
rect 4340 14662 4362 14714
rect 4362 14662 4374 14714
rect 4374 14662 4396 14714
rect 4420 14662 4426 14714
rect 4426 14662 4438 14714
rect 4438 14662 4476 14714
rect 4500 14662 4502 14714
rect 4502 14662 4554 14714
rect 4554 14662 4556 14714
rect 4180 14660 4236 14662
rect 4260 14660 4316 14662
rect 4340 14660 4396 14662
rect 4420 14660 4476 14662
rect 4500 14660 4556 14662
rect 4920 16346 4976 16348
rect 5000 16346 5056 16348
rect 5080 16346 5136 16348
rect 5160 16346 5216 16348
rect 5240 16346 5296 16348
rect 4920 16294 4922 16346
rect 4922 16294 4974 16346
rect 4974 16294 4976 16346
rect 5000 16294 5038 16346
rect 5038 16294 5050 16346
rect 5050 16294 5056 16346
rect 5080 16294 5102 16346
rect 5102 16294 5114 16346
rect 5114 16294 5136 16346
rect 5160 16294 5166 16346
rect 5166 16294 5178 16346
rect 5178 16294 5216 16346
rect 5240 16294 5242 16346
rect 5242 16294 5294 16346
rect 5294 16294 5296 16346
rect 4920 16292 4976 16294
rect 5000 16292 5056 16294
rect 5080 16292 5136 16294
rect 5160 16292 5216 16294
rect 5240 16292 5296 16294
rect 4920 15258 4976 15260
rect 5000 15258 5056 15260
rect 5080 15258 5136 15260
rect 5160 15258 5216 15260
rect 5240 15258 5296 15260
rect 4920 15206 4922 15258
rect 4922 15206 4974 15258
rect 4974 15206 4976 15258
rect 5000 15206 5038 15258
rect 5038 15206 5050 15258
rect 5050 15206 5056 15258
rect 5080 15206 5102 15258
rect 5102 15206 5114 15258
rect 5114 15206 5136 15258
rect 5160 15206 5166 15258
rect 5166 15206 5178 15258
rect 5178 15206 5216 15258
rect 5240 15206 5242 15258
rect 5242 15206 5294 15258
rect 5294 15206 5296 15258
rect 4920 15204 4976 15206
rect 5000 15204 5056 15206
rect 5080 15204 5136 15206
rect 5160 15204 5216 15206
rect 5240 15204 5296 15206
rect 4180 13626 4236 13628
rect 4260 13626 4316 13628
rect 4340 13626 4396 13628
rect 4420 13626 4476 13628
rect 4500 13626 4556 13628
rect 4180 13574 4182 13626
rect 4182 13574 4234 13626
rect 4234 13574 4236 13626
rect 4260 13574 4298 13626
rect 4298 13574 4310 13626
rect 4310 13574 4316 13626
rect 4340 13574 4362 13626
rect 4362 13574 4374 13626
rect 4374 13574 4396 13626
rect 4420 13574 4426 13626
rect 4426 13574 4438 13626
rect 4438 13574 4476 13626
rect 4500 13574 4502 13626
rect 4502 13574 4554 13626
rect 4554 13574 4556 13626
rect 4180 13572 4236 13574
rect 4260 13572 4316 13574
rect 4340 13572 4396 13574
rect 4420 13572 4476 13574
rect 4500 13572 4556 13574
rect 4180 12538 4236 12540
rect 4260 12538 4316 12540
rect 4340 12538 4396 12540
rect 4420 12538 4476 12540
rect 4500 12538 4556 12540
rect 4180 12486 4182 12538
rect 4182 12486 4234 12538
rect 4234 12486 4236 12538
rect 4260 12486 4298 12538
rect 4298 12486 4310 12538
rect 4310 12486 4316 12538
rect 4340 12486 4362 12538
rect 4362 12486 4374 12538
rect 4374 12486 4396 12538
rect 4420 12486 4426 12538
rect 4426 12486 4438 12538
rect 4438 12486 4476 12538
rect 4500 12486 4502 12538
rect 4502 12486 4554 12538
rect 4554 12486 4556 12538
rect 4180 12484 4236 12486
rect 4260 12484 4316 12486
rect 4340 12484 4396 12486
rect 4420 12484 4476 12486
rect 4500 12484 4556 12486
rect 4920 14170 4976 14172
rect 5000 14170 5056 14172
rect 5080 14170 5136 14172
rect 5160 14170 5216 14172
rect 5240 14170 5296 14172
rect 4920 14118 4922 14170
rect 4922 14118 4974 14170
rect 4974 14118 4976 14170
rect 5000 14118 5038 14170
rect 5038 14118 5050 14170
rect 5050 14118 5056 14170
rect 5080 14118 5102 14170
rect 5102 14118 5114 14170
rect 5114 14118 5136 14170
rect 5160 14118 5166 14170
rect 5166 14118 5178 14170
rect 5178 14118 5216 14170
rect 5240 14118 5242 14170
rect 5242 14118 5294 14170
rect 5294 14118 5296 14170
rect 4920 14116 4976 14118
rect 5000 14116 5056 14118
rect 5080 14116 5136 14118
rect 5160 14116 5216 14118
rect 5240 14116 5296 14118
rect 4920 13082 4976 13084
rect 5000 13082 5056 13084
rect 5080 13082 5136 13084
rect 5160 13082 5216 13084
rect 5240 13082 5296 13084
rect 4920 13030 4922 13082
rect 4922 13030 4974 13082
rect 4974 13030 4976 13082
rect 5000 13030 5038 13082
rect 5038 13030 5050 13082
rect 5050 13030 5056 13082
rect 5080 13030 5102 13082
rect 5102 13030 5114 13082
rect 5114 13030 5136 13082
rect 5160 13030 5166 13082
rect 5166 13030 5178 13082
rect 5178 13030 5216 13082
rect 5240 13030 5242 13082
rect 5242 13030 5294 13082
rect 5294 13030 5296 13082
rect 4920 13028 4976 13030
rect 5000 13028 5056 13030
rect 5080 13028 5136 13030
rect 5160 13028 5216 13030
rect 5240 13028 5296 13030
rect 4180 11450 4236 11452
rect 4260 11450 4316 11452
rect 4340 11450 4396 11452
rect 4420 11450 4476 11452
rect 4500 11450 4556 11452
rect 4180 11398 4182 11450
rect 4182 11398 4234 11450
rect 4234 11398 4236 11450
rect 4260 11398 4298 11450
rect 4298 11398 4310 11450
rect 4310 11398 4316 11450
rect 4340 11398 4362 11450
rect 4362 11398 4374 11450
rect 4374 11398 4396 11450
rect 4420 11398 4426 11450
rect 4426 11398 4438 11450
rect 4438 11398 4476 11450
rect 4500 11398 4502 11450
rect 4502 11398 4554 11450
rect 4554 11398 4556 11450
rect 4180 11396 4236 11398
rect 4260 11396 4316 11398
rect 4340 11396 4396 11398
rect 4420 11396 4476 11398
rect 4500 11396 4556 11398
rect 4920 11994 4976 11996
rect 5000 11994 5056 11996
rect 5080 11994 5136 11996
rect 5160 11994 5216 11996
rect 5240 11994 5296 11996
rect 4920 11942 4922 11994
rect 4922 11942 4974 11994
rect 4974 11942 4976 11994
rect 5000 11942 5038 11994
rect 5038 11942 5050 11994
rect 5050 11942 5056 11994
rect 5080 11942 5102 11994
rect 5102 11942 5114 11994
rect 5114 11942 5136 11994
rect 5160 11942 5166 11994
rect 5166 11942 5178 11994
rect 5178 11942 5216 11994
rect 5240 11942 5242 11994
rect 5242 11942 5294 11994
rect 5294 11942 5296 11994
rect 4920 11940 4976 11942
rect 5000 11940 5056 11942
rect 5080 11940 5136 11942
rect 5160 11940 5216 11942
rect 5240 11940 5296 11942
rect 10920 30490 10976 30492
rect 11000 30490 11056 30492
rect 11080 30490 11136 30492
rect 11160 30490 11216 30492
rect 11240 30490 11296 30492
rect 10920 30438 10922 30490
rect 10922 30438 10974 30490
rect 10974 30438 10976 30490
rect 11000 30438 11038 30490
rect 11038 30438 11050 30490
rect 11050 30438 11056 30490
rect 11080 30438 11102 30490
rect 11102 30438 11114 30490
rect 11114 30438 11136 30490
rect 11160 30438 11166 30490
rect 11166 30438 11178 30490
rect 11178 30438 11216 30490
rect 11240 30438 11242 30490
rect 11242 30438 11294 30490
rect 11294 30438 11296 30490
rect 10920 30436 10976 30438
rect 11000 30436 11056 30438
rect 11080 30436 11136 30438
rect 11160 30436 11216 30438
rect 11240 30436 11296 30438
rect 10920 29402 10976 29404
rect 11000 29402 11056 29404
rect 11080 29402 11136 29404
rect 11160 29402 11216 29404
rect 11240 29402 11296 29404
rect 10920 29350 10922 29402
rect 10922 29350 10974 29402
rect 10974 29350 10976 29402
rect 11000 29350 11038 29402
rect 11038 29350 11050 29402
rect 11050 29350 11056 29402
rect 11080 29350 11102 29402
rect 11102 29350 11114 29402
rect 11114 29350 11136 29402
rect 11160 29350 11166 29402
rect 11166 29350 11178 29402
rect 11178 29350 11216 29402
rect 11240 29350 11242 29402
rect 11242 29350 11294 29402
rect 11294 29350 11296 29402
rect 10920 29348 10976 29350
rect 11000 29348 11056 29350
rect 11080 29348 11136 29350
rect 11160 29348 11216 29350
rect 11240 29348 11296 29350
rect 9218 26968 9274 27024
rect 8206 21548 8262 21584
rect 8206 21528 8208 21548
rect 8208 21528 8260 21548
rect 8260 21528 8262 21548
rect 10180 27770 10236 27772
rect 10260 27770 10316 27772
rect 10340 27770 10396 27772
rect 10420 27770 10476 27772
rect 10500 27770 10556 27772
rect 10180 27718 10182 27770
rect 10182 27718 10234 27770
rect 10234 27718 10236 27770
rect 10260 27718 10298 27770
rect 10298 27718 10310 27770
rect 10310 27718 10316 27770
rect 10340 27718 10362 27770
rect 10362 27718 10374 27770
rect 10374 27718 10396 27770
rect 10420 27718 10426 27770
rect 10426 27718 10438 27770
rect 10438 27718 10476 27770
rect 10500 27718 10502 27770
rect 10502 27718 10554 27770
rect 10554 27718 10556 27770
rect 10180 27716 10236 27718
rect 10260 27716 10316 27718
rect 10340 27716 10396 27718
rect 10420 27716 10476 27718
rect 10500 27716 10556 27718
rect 10180 26682 10236 26684
rect 10260 26682 10316 26684
rect 10340 26682 10396 26684
rect 10420 26682 10476 26684
rect 10500 26682 10556 26684
rect 10180 26630 10182 26682
rect 10182 26630 10234 26682
rect 10234 26630 10236 26682
rect 10260 26630 10298 26682
rect 10298 26630 10310 26682
rect 10310 26630 10316 26682
rect 10340 26630 10362 26682
rect 10362 26630 10374 26682
rect 10374 26630 10396 26682
rect 10420 26630 10426 26682
rect 10426 26630 10438 26682
rect 10438 26630 10476 26682
rect 10500 26630 10502 26682
rect 10502 26630 10554 26682
rect 10554 26630 10556 26682
rect 10180 26628 10236 26630
rect 10260 26628 10316 26630
rect 10340 26628 10396 26630
rect 10420 26628 10476 26630
rect 10500 26628 10556 26630
rect 10180 25594 10236 25596
rect 10260 25594 10316 25596
rect 10340 25594 10396 25596
rect 10420 25594 10476 25596
rect 10500 25594 10556 25596
rect 10180 25542 10182 25594
rect 10182 25542 10234 25594
rect 10234 25542 10236 25594
rect 10260 25542 10298 25594
rect 10298 25542 10310 25594
rect 10310 25542 10316 25594
rect 10340 25542 10362 25594
rect 10362 25542 10374 25594
rect 10374 25542 10396 25594
rect 10420 25542 10426 25594
rect 10426 25542 10438 25594
rect 10438 25542 10476 25594
rect 10500 25542 10502 25594
rect 10502 25542 10554 25594
rect 10554 25542 10556 25594
rect 10180 25540 10236 25542
rect 10260 25540 10316 25542
rect 10340 25540 10396 25542
rect 10420 25540 10476 25542
rect 10500 25540 10556 25542
rect 10920 28314 10976 28316
rect 11000 28314 11056 28316
rect 11080 28314 11136 28316
rect 11160 28314 11216 28316
rect 11240 28314 11296 28316
rect 10920 28262 10922 28314
rect 10922 28262 10974 28314
rect 10974 28262 10976 28314
rect 11000 28262 11038 28314
rect 11038 28262 11050 28314
rect 11050 28262 11056 28314
rect 11080 28262 11102 28314
rect 11102 28262 11114 28314
rect 11114 28262 11136 28314
rect 11160 28262 11166 28314
rect 11166 28262 11178 28314
rect 11178 28262 11216 28314
rect 11240 28262 11242 28314
rect 11242 28262 11294 28314
rect 11294 28262 11296 28314
rect 10920 28260 10976 28262
rect 11000 28260 11056 28262
rect 11080 28260 11136 28262
rect 11160 28260 11216 28262
rect 11240 28260 11296 28262
rect 10920 27226 10976 27228
rect 11000 27226 11056 27228
rect 11080 27226 11136 27228
rect 11160 27226 11216 27228
rect 11240 27226 11296 27228
rect 10920 27174 10922 27226
rect 10922 27174 10974 27226
rect 10974 27174 10976 27226
rect 11000 27174 11038 27226
rect 11038 27174 11050 27226
rect 11050 27174 11056 27226
rect 11080 27174 11102 27226
rect 11102 27174 11114 27226
rect 11114 27174 11136 27226
rect 11160 27174 11166 27226
rect 11166 27174 11178 27226
rect 11178 27174 11216 27226
rect 11240 27174 11242 27226
rect 11242 27174 11294 27226
rect 11294 27174 11296 27226
rect 10920 27172 10976 27174
rect 11000 27172 11056 27174
rect 11080 27172 11136 27174
rect 11160 27172 11216 27174
rect 11240 27172 11296 27174
rect 10920 26138 10976 26140
rect 11000 26138 11056 26140
rect 11080 26138 11136 26140
rect 11160 26138 11216 26140
rect 11240 26138 11296 26140
rect 10920 26086 10922 26138
rect 10922 26086 10974 26138
rect 10974 26086 10976 26138
rect 11000 26086 11038 26138
rect 11038 26086 11050 26138
rect 11050 26086 11056 26138
rect 11080 26086 11102 26138
rect 11102 26086 11114 26138
rect 11114 26086 11136 26138
rect 11160 26086 11166 26138
rect 11166 26086 11178 26138
rect 11178 26086 11216 26138
rect 11240 26086 11242 26138
rect 11242 26086 11294 26138
rect 11294 26086 11296 26138
rect 10920 26084 10976 26086
rect 11000 26084 11056 26086
rect 11080 26084 11136 26086
rect 11160 26084 11216 26086
rect 11240 26084 11296 26086
rect 10690 24676 10746 24712
rect 10690 24656 10692 24676
rect 10692 24656 10744 24676
rect 10744 24656 10746 24676
rect 10180 24506 10236 24508
rect 10260 24506 10316 24508
rect 10340 24506 10396 24508
rect 10420 24506 10476 24508
rect 10500 24506 10556 24508
rect 10180 24454 10182 24506
rect 10182 24454 10234 24506
rect 10234 24454 10236 24506
rect 10260 24454 10298 24506
rect 10298 24454 10310 24506
rect 10310 24454 10316 24506
rect 10340 24454 10362 24506
rect 10362 24454 10374 24506
rect 10374 24454 10396 24506
rect 10420 24454 10426 24506
rect 10426 24454 10438 24506
rect 10438 24454 10476 24506
rect 10500 24454 10502 24506
rect 10502 24454 10554 24506
rect 10554 24454 10556 24506
rect 10180 24452 10236 24454
rect 10260 24452 10316 24454
rect 10340 24452 10396 24454
rect 10420 24452 10476 24454
rect 10500 24452 10556 24454
rect 10180 23418 10236 23420
rect 10260 23418 10316 23420
rect 10340 23418 10396 23420
rect 10420 23418 10476 23420
rect 10500 23418 10556 23420
rect 10180 23366 10182 23418
rect 10182 23366 10234 23418
rect 10234 23366 10236 23418
rect 10260 23366 10298 23418
rect 10298 23366 10310 23418
rect 10310 23366 10316 23418
rect 10340 23366 10362 23418
rect 10362 23366 10374 23418
rect 10374 23366 10396 23418
rect 10420 23366 10426 23418
rect 10426 23366 10438 23418
rect 10438 23366 10476 23418
rect 10500 23366 10502 23418
rect 10502 23366 10554 23418
rect 10554 23366 10556 23418
rect 10180 23364 10236 23366
rect 10260 23364 10316 23366
rect 10340 23364 10396 23366
rect 10420 23364 10476 23366
rect 10500 23364 10556 23366
rect 10180 22330 10236 22332
rect 10260 22330 10316 22332
rect 10340 22330 10396 22332
rect 10420 22330 10476 22332
rect 10500 22330 10556 22332
rect 10180 22278 10182 22330
rect 10182 22278 10234 22330
rect 10234 22278 10236 22330
rect 10260 22278 10298 22330
rect 10298 22278 10310 22330
rect 10310 22278 10316 22330
rect 10340 22278 10362 22330
rect 10362 22278 10374 22330
rect 10374 22278 10396 22330
rect 10420 22278 10426 22330
rect 10426 22278 10438 22330
rect 10438 22278 10476 22330
rect 10500 22278 10502 22330
rect 10502 22278 10554 22330
rect 10554 22278 10556 22330
rect 10180 22276 10236 22278
rect 10260 22276 10316 22278
rect 10340 22276 10396 22278
rect 10420 22276 10476 22278
rect 10500 22276 10556 22278
rect 10180 21242 10236 21244
rect 10260 21242 10316 21244
rect 10340 21242 10396 21244
rect 10420 21242 10476 21244
rect 10500 21242 10556 21244
rect 10180 21190 10182 21242
rect 10182 21190 10234 21242
rect 10234 21190 10236 21242
rect 10260 21190 10298 21242
rect 10298 21190 10310 21242
rect 10310 21190 10316 21242
rect 10340 21190 10362 21242
rect 10362 21190 10374 21242
rect 10374 21190 10396 21242
rect 10420 21190 10426 21242
rect 10426 21190 10438 21242
rect 10438 21190 10476 21242
rect 10500 21190 10502 21242
rect 10502 21190 10554 21242
rect 10554 21190 10556 21242
rect 10180 21188 10236 21190
rect 10260 21188 10316 21190
rect 10340 21188 10396 21190
rect 10420 21188 10476 21190
rect 10500 21188 10556 21190
rect 10920 25050 10976 25052
rect 11000 25050 11056 25052
rect 11080 25050 11136 25052
rect 11160 25050 11216 25052
rect 11240 25050 11296 25052
rect 10920 24998 10922 25050
rect 10922 24998 10974 25050
rect 10974 24998 10976 25050
rect 11000 24998 11038 25050
rect 11038 24998 11050 25050
rect 11050 24998 11056 25050
rect 11080 24998 11102 25050
rect 11102 24998 11114 25050
rect 11114 24998 11136 25050
rect 11160 24998 11166 25050
rect 11166 24998 11178 25050
rect 11178 24998 11216 25050
rect 11240 24998 11242 25050
rect 11242 24998 11294 25050
rect 11294 24998 11296 25050
rect 10920 24996 10976 24998
rect 11000 24996 11056 24998
rect 11080 24996 11136 24998
rect 11160 24996 11216 24998
rect 11240 24996 11296 24998
rect 10920 23962 10976 23964
rect 11000 23962 11056 23964
rect 11080 23962 11136 23964
rect 11160 23962 11216 23964
rect 11240 23962 11296 23964
rect 10920 23910 10922 23962
rect 10922 23910 10974 23962
rect 10974 23910 10976 23962
rect 11000 23910 11038 23962
rect 11038 23910 11050 23962
rect 11050 23910 11056 23962
rect 11080 23910 11102 23962
rect 11102 23910 11114 23962
rect 11114 23910 11136 23962
rect 11160 23910 11166 23962
rect 11166 23910 11178 23962
rect 11178 23910 11216 23962
rect 11240 23910 11242 23962
rect 11242 23910 11294 23962
rect 11294 23910 11296 23962
rect 10920 23908 10976 23910
rect 11000 23908 11056 23910
rect 11080 23908 11136 23910
rect 11160 23908 11216 23910
rect 11240 23908 11296 23910
rect 10920 22874 10976 22876
rect 11000 22874 11056 22876
rect 11080 22874 11136 22876
rect 11160 22874 11216 22876
rect 11240 22874 11296 22876
rect 10920 22822 10922 22874
rect 10922 22822 10974 22874
rect 10974 22822 10976 22874
rect 11000 22822 11038 22874
rect 11038 22822 11050 22874
rect 11050 22822 11056 22874
rect 11080 22822 11102 22874
rect 11102 22822 11114 22874
rect 11114 22822 11136 22874
rect 11160 22822 11166 22874
rect 11166 22822 11178 22874
rect 11178 22822 11216 22874
rect 11240 22822 11242 22874
rect 11242 22822 11294 22874
rect 11294 22822 11296 22874
rect 10920 22820 10976 22822
rect 11000 22820 11056 22822
rect 11080 22820 11136 22822
rect 11160 22820 11216 22822
rect 11240 22820 11296 22822
rect 10920 21786 10976 21788
rect 11000 21786 11056 21788
rect 11080 21786 11136 21788
rect 11160 21786 11216 21788
rect 11240 21786 11296 21788
rect 10920 21734 10922 21786
rect 10922 21734 10974 21786
rect 10974 21734 10976 21786
rect 11000 21734 11038 21786
rect 11038 21734 11050 21786
rect 11050 21734 11056 21786
rect 11080 21734 11102 21786
rect 11102 21734 11114 21786
rect 11114 21734 11136 21786
rect 11160 21734 11166 21786
rect 11166 21734 11178 21786
rect 11178 21734 11216 21786
rect 11240 21734 11242 21786
rect 11242 21734 11294 21786
rect 11294 21734 11296 21786
rect 10920 21732 10976 21734
rect 11000 21732 11056 21734
rect 11080 21732 11136 21734
rect 11160 21732 11216 21734
rect 11240 21732 11296 21734
rect 11334 21528 11390 21584
rect 4920 10906 4976 10908
rect 5000 10906 5056 10908
rect 5080 10906 5136 10908
rect 5160 10906 5216 10908
rect 5240 10906 5296 10908
rect 4920 10854 4922 10906
rect 4922 10854 4974 10906
rect 4974 10854 4976 10906
rect 5000 10854 5038 10906
rect 5038 10854 5050 10906
rect 5050 10854 5056 10906
rect 5080 10854 5102 10906
rect 5102 10854 5114 10906
rect 5114 10854 5136 10906
rect 5160 10854 5166 10906
rect 5166 10854 5178 10906
rect 5178 10854 5216 10906
rect 5240 10854 5242 10906
rect 5242 10854 5294 10906
rect 5294 10854 5296 10906
rect 4920 10852 4976 10854
rect 5000 10852 5056 10854
rect 5080 10852 5136 10854
rect 5160 10852 5216 10854
rect 5240 10852 5296 10854
rect 4180 10362 4236 10364
rect 4260 10362 4316 10364
rect 4340 10362 4396 10364
rect 4420 10362 4476 10364
rect 4500 10362 4556 10364
rect 4180 10310 4182 10362
rect 4182 10310 4234 10362
rect 4234 10310 4236 10362
rect 4260 10310 4298 10362
rect 4298 10310 4310 10362
rect 4310 10310 4316 10362
rect 4340 10310 4362 10362
rect 4362 10310 4374 10362
rect 4374 10310 4396 10362
rect 4420 10310 4426 10362
rect 4426 10310 4438 10362
rect 4438 10310 4476 10362
rect 4500 10310 4502 10362
rect 4502 10310 4554 10362
rect 4554 10310 4556 10362
rect 4180 10308 4236 10310
rect 4260 10308 4316 10310
rect 4340 10308 4396 10310
rect 4420 10308 4476 10310
rect 4500 10308 4556 10310
rect 4180 9274 4236 9276
rect 4260 9274 4316 9276
rect 4340 9274 4396 9276
rect 4420 9274 4476 9276
rect 4500 9274 4556 9276
rect 4180 9222 4182 9274
rect 4182 9222 4234 9274
rect 4234 9222 4236 9274
rect 4260 9222 4298 9274
rect 4298 9222 4310 9274
rect 4310 9222 4316 9274
rect 4340 9222 4362 9274
rect 4362 9222 4374 9274
rect 4374 9222 4396 9274
rect 4420 9222 4426 9274
rect 4426 9222 4438 9274
rect 4438 9222 4476 9274
rect 4500 9222 4502 9274
rect 4502 9222 4554 9274
rect 4554 9222 4556 9274
rect 4180 9220 4236 9222
rect 4260 9220 4316 9222
rect 4340 9220 4396 9222
rect 4420 9220 4476 9222
rect 4500 9220 4556 9222
rect 4180 8186 4236 8188
rect 4260 8186 4316 8188
rect 4340 8186 4396 8188
rect 4420 8186 4476 8188
rect 4500 8186 4556 8188
rect 4180 8134 4182 8186
rect 4182 8134 4234 8186
rect 4234 8134 4236 8186
rect 4260 8134 4298 8186
rect 4298 8134 4310 8186
rect 4310 8134 4316 8186
rect 4340 8134 4362 8186
rect 4362 8134 4374 8186
rect 4374 8134 4396 8186
rect 4420 8134 4426 8186
rect 4426 8134 4438 8186
rect 4438 8134 4476 8186
rect 4500 8134 4502 8186
rect 4502 8134 4554 8186
rect 4554 8134 4556 8186
rect 4180 8132 4236 8134
rect 4260 8132 4316 8134
rect 4340 8132 4396 8134
rect 4420 8132 4476 8134
rect 4500 8132 4556 8134
rect 4180 7098 4236 7100
rect 4260 7098 4316 7100
rect 4340 7098 4396 7100
rect 4420 7098 4476 7100
rect 4500 7098 4556 7100
rect 4180 7046 4182 7098
rect 4182 7046 4234 7098
rect 4234 7046 4236 7098
rect 4260 7046 4298 7098
rect 4298 7046 4310 7098
rect 4310 7046 4316 7098
rect 4340 7046 4362 7098
rect 4362 7046 4374 7098
rect 4374 7046 4396 7098
rect 4420 7046 4426 7098
rect 4426 7046 4438 7098
rect 4438 7046 4476 7098
rect 4500 7046 4502 7098
rect 4502 7046 4554 7098
rect 4554 7046 4556 7098
rect 4180 7044 4236 7046
rect 4260 7044 4316 7046
rect 4340 7044 4396 7046
rect 4420 7044 4476 7046
rect 4500 7044 4556 7046
rect 4920 9818 4976 9820
rect 5000 9818 5056 9820
rect 5080 9818 5136 9820
rect 5160 9818 5216 9820
rect 5240 9818 5296 9820
rect 4920 9766 4922 9818
rect 4922 9766 4974 9818
rect 4974 9766 4976 9818
rect 5000 9766 5038 9818
rect 5038 9766 5050 9818
rect 5050 9766 5056 9818
rect 5080 9766 5102 9818
rect 5102 9766 5114 9818
rect 5114 9766 5136 9818
rect 5160 9766 5166 9818
rect 5166 9766 5178 9818
rect 5178 9766 5216 9818
rect 5240 9766 5242 9818
rect 5242 9766 5294 9818
rect 5294 9766 5296 9818
rect 4920 9764 4976 9766
rect 5000 9764 5056 9766
rect 5080 9764 5136 9766
rect 5160 9764 5216 9766
rect 5240 9764 5296 9766
rect 4920 8730 4976 8732
rect 5000 8730 5056 8732
rect 5080 8730 5136 8732
rect 5160 8730 5216 8732
rect 5240 8730 5296 8732
rect 4920 8678 4922 8730
rect 4922 8678 4974 8730
rect 4974 8678 4976 8730
rect 5000 8678 5038 8730
rect 5038 8678 5050 8730
rect 5050 8678 5056 8730
rect 5080 8678 5102 8730
rect 5102 8678 5114 8730
rect 5114 8678 5136 8730
rect 5160 8678 5166 8730
rect 5166 8678 5178 8730
rect 5178 8678 5216 8730
rect 5240 8678 5242 8730
rect 5242 8678 5294 8730
rect 5294 8678 5296 8730
rect 4920 8676 4976 8678
rect 5000 8676 5056 8678
rect 5080 8676 5136 8678
rect 5160 8676 5216 8678
rect 5240 8676 5296 8678
rect 4920 7642 4976 7644
rect 5000 7642 5056 7644
rect 5080 7642 5136 7644
rect 5160 7642 5216 7644
rect 5240 7642 5296 7644
rect 4920 7590 4922 7642
rect 4922 7590 4974 7642
rect 4974 7590 4976 7642
rect 5000 7590 5038 7642
rect 5038 7590 5050 7642
rect 5050 7590 5056 7642
rect 5080 7590 5102 7642
rect 5102 7590 5114 7642
rect 5114 7590 5136 7642
rect 5160 7590 5166 7642
rect 5166 7590 5178 7642
rect 5178 7590 5216 7642
rect 5240 7590 5242 7642
rect 5242 7590 5294 7642
rect 5294 7590 5296 7642
rect 4920 7588 4976 7590
rect 5000 7588 5056 7590
rect 5080 7588 5136 7590
rect 5160 7588 5216 7590
rect 5240 7588 5296 7590
rect 4920 6554 4976 6556
rect 5000 6554 5056 6556
rect 5080 6554 5136 6556
rect 5160 6554 5216 6556
rect 5240 6554 5296 6556
rect 4920 6502 4922 6554
rect 4922 6502 4974 6554
rect 4974 6502 4976 6554
rect 5000 6502 5038 6554
rect 5038 6502 5050 6554
rect 5050 6502 5056 6554
rect 5080 6502 5102 6554
rect 5102 6502 5114 6554
rect 5114 6502 5136 6554
rect 5160 6502 5166 6554
rect 5166 6502 5178 6554
rect 5178 6502 5216 6554
rect 5240 6502 5242 6554
rect 5242 6502 5294 6554
rect 5294 6502 5296 6554
rect 4920 6500 4976 6502
rect 5000 6500 5056 6502
rect 5080 6500 5136 6502
rect 5160 6500 5216 6502
rect 5240 6500 5296 6502
rect 938 6160 994 6216
rect 4180 6010 4236 6012
rect 4260 6010 4316 6012
rect 4340 6010 4396 6012
rect 4420 6010 4476 6012
rect 4500 6010 4556 6012
rect 4180 5958 4182 6010
rect 4182 5958 4234 6010
rect 4234 5958 4236 6010
rect 4260 5958 4298 6010
rect 4298 5958 4310 6010
rect 4310 5958 4316 6010
rect 4340 5958 4362 6010
rect 4362 5958 4374 6010
rect 4374 5958 4396 6010
rect 4420 5958 4426 6010
rect 4426 5958 4438 6010
rect 4438 5958 4476 6010
rect 4500 5958 4502 6010
rect 4502 5958 4554 6010
rect 4554 5958 4556 6010
rect 4180 5956 4236 5958
rect 4260 5956 4316 5958
rect 4340 5956 4396 5958
rect 4420 5956 4476 5958
rect 4500 5956 4556 5958
rect 10180 20154 10236 20156
rect 10260 20154 10316 20156
rect 10340 20154 10396 20156
rect 10420 20154 10476 20156
rect 10500 20154 10556 20156
rect 10180 20102 10182 20154
rect 10182 20102 10234 20154
rect 10234 20102 10236 20154
rect 10260 20102 10298 20154
rect 10298 20102 10310 20154
rect 10310 20102 10316 20154
rect 10340 20102 10362 20154
rect 10362 20102 10374 20154
rect 10374 20102 10396 20154
rect 10420 20102 10426 20154
rect 10426 20102 10438 20154
rect 10438 20102 10476 20154
rect 10500 20102 10502 20154
rect 10502 20102 10554 20154
rect 10554 20102 10556 20154
rect 10180 20100 10236 20102
rect 10260 20100 10316 20102
rect 10340 20100 10396 20102
rect 10420 20100 10476 20102
rect 10500 20100 10556 20102
rect 10180 19066 10236 19068
rect 10260 19066 10316 19068
rect 10340 19066 10396 19068
rect 10420 19066 10476 19068
rect 10500 19066 10556 19068
rect 10180 19014 10182 19066
rect 10182 19014 10234 19066
rect 10234 19014 10236 19066
rect 10260 19014 10298 19066
rect 10298 19014 10310 19066
rect 10310 19014 10316 19066
rect 10340 19014 10362 19066
rect 10362 19014 10374 19066
rect 10374 19014 10396 19066
rect 10420 19014 10426 19066
rect 10426 19014 10438 19066
rect 10438 19014 10476 19066
rect 10500 19014 10502 19066
rect 10502 19014 10554 19066
rect 10554 19014 10556 19066
rect 10180 19012 10236 19014
rect 10260 19012 10316 19014
rect 10340 19012 10396 19014
rect 10420 19012 10476 19014
rect 10500 19012 10556 19014
rect 10920 20698 10976 20700
rect 11000 20698 11056 20700
rect 11080 20698 11136 20700
rect 11160 20698 11216 20700
rect 11240 20698 11296 20700
rect 10920 20646 10922 20698
rect 10922 20646 10974 20698
rect 10974 20646 10976 20698
rect 11000 20646 11038 20698
rect 11038 20646 11050 20698
rect 11050 20646 11056 20698
rect 11080 20646 11102 20698
rect 11102 20646 11114 20698
rect 11114 20646 11136 20698
rect 11160 20646 11166 20698
rect 11166 20646 11178 20698
rect 11178 20646 11216 20698
rect 11240 20646 11242 20698
rect 11242 20646 11294 20698
rect 11294 20646 11296 20698
rect 10920 20644 10976 20646
rect 11000 20644 11056 20646
rect 11080 20644 11136 20646
rect 11160 20644 11216 20646
rect 11240 20644 11296 20646
rect 4920 5466 4976 5468
rect 5000 5466 5056 5468
rect 5080 5466 5136 5468
rect 5160 5466 5216 5468
rect 5240 5466 5296 5468
rect 4920 5414 4922 5466
rect 4922 5414 4974 5466
rect 4974 5414 4976 5466
rect 5000 5414 5038 5466
rect 5038 5414 5050 5466
rect 5050 5414 5056 5466
rect 5080 5414 5102 5466
rect 5102 5414 5114 5466
rect 5114 5414 5136 5466
rect 5160 5414 5166 5466
rect 5166 5414 5178 5466
rect 5178 5414 5216 5466
rect 5240 5414 5242 5466
rect 5242 5414 5294 5466
rect 5294 5414 5296 5466
rect 4920 5412 4976 5414
rect 5000 5412 5056 5414
rect 5080 5412 5136 5414
rect 5160 5412 5216 5414
rect 5240 5412 5296 5414
rect 4180 4922 4236 4924
rect 4260 4922 4316 4924
rect 4340 4922 4396 4924
rect 4420 4922 4476 4924
rect 4500 4922 4556 4924
rect 4180 4870 4182 4922
rect 4182 4870 4234 4922
rect 4234 4870 4236 4922
rect 4260 4870 4298 4922
rect 4298 4870 4310 4922
rect 4310 4870 4316 4922
rect 4340 4870 4362 4922
rect 4362 4870 4374 4922
rect 4374 4870 4396 4922
rect 4420 4870 4426 4922
rect 4426 4870 4438 4922
rect 4438 4870 4476 4922
rect 4500 4870 4502 4922
rect 4502 4870 4554 4922
rect 4554 4870 4556 4922
rect 4180 4868 4236 4870
rect 4260 4868 4316 4870
rect 4340 4868 4396 4870
rect 4420 4868 4476 4870
rect 4500 4868 4556 4870
rect 4920 4378 4976 4380
rect 5000 4378 5056 4380
rect 5080 4378 5136 4380
rect 5160 4378 5216 4380
rect 5240 4378 5296 4380
rect 4920 4326 4922 4378
rect 4922 4326 4974 4378
rect 4974 4326 4976 4378
rect 5000 4326 5038 4378
rect 5038 4326 5050 4378
rect 5050 4326 5056 4378
rect 5080 4326 5102 4378
rect 5102 4326 5114 4378
rect 5114 4326 5136 4378
rect 5160 4326 5166 4378
rect 5166 4326 5178 4378
rect 5178 4326 5216 4378
rect 5240 4326 5242 4378
rect 5242 4326 5294 4378
rect 5294 4326 5296 4378
rect 4920 4324 4976 4326
rect 5000 4324 5056 4326
rect 5080 4324 5136 4326
rect 5160 4324 5216 4326
rect 5240 4324 5296 4326
rect 10180 17978 10236 17980
rect 10260 17978 10316 17980
rect 10340 17978 10396 17980
rect 10420 17978 10476 17980
rect 10500 17978 10556 17980
rect 10180 17926 10182 17978
rect 10182 17926 10234 17978
rect 10234 17926 10236 17978
rect 10260 17926 10298 17978
rect 10298 17926 10310 17978
rect 10310 17926 10316 17978
rect 10340 17926 10362 17978
rect 10362 17926 10374 17978
rect 10374 17926 10396 17978
rect 10420 17926 10426 17978
rect 10426 17926 10438 17978
rect 10438 17926 10476 17978
rect 10500 17926 10502 17978
rect 10502 17926 10554 17978
rect 10554 17926 10556 17978
rect 10180 17924 10236 17926
rect 10260 17924 10316 17926
rect 10340 17924 10396 17926
rect 10420 17924 10476 17926
rect 10500 17924 10556 17926
rect 10180 16890 10236 16892
rect 10260 16890 10316 16892
rect 10340 16890 10396 16892
rect 10420 16890 10476 16892
rect 10500 16890 10556 16892
rect 10180 16838 10182 16890
rect 10182 16838 10234 16890
rect 10234 16838 10236 16890
rect 10260 16838 10298 16890
rect 10298 16838 10310 16890
rect 10310 16838 10316 16890
rect 10340 16838 10362 16890
rect 10362 16838 10374 16890
rect 10374 16838 10396 16890
rect 10420 16838 10426 16890
rect 10426 16838 10438 16890
rect 10438 16838 10476 16890
rect 10500 16838 10502 16890
rect 10502 16838 10554 16890
rect 10554 16838 10556 16890
rect 10180 16836 10236 16838
rect 10260 16836 10316 16838
rect 10340 16836 10396 16838
rect 10420 16836 10476 16838
rect 10500 16836 10556 16838
rect 10180 15802 10236 15804
rect 10260 15802 10316 15804
rect 10340 15802 10396 15804
rect 10420 15802 10476 15804
rect 10500 15802 10556 15804
rect 10180 15750 10182 15802
rect 10182 15750 10234 15802
rect 10234 15750 10236 15802
rect 10260 15750 10298 15802
rect 10298 15750 10310 15802
rect 10310 15750 10316 15802
rect 10340 15750 10362 15802
rect 10362 15750 10374 15802
rect 10374 15750 10396 15802
rect 10420 15750 10426 15802
rect 10426 15750 10438 15802
rect 10438 15750 10476 15802
rect 10500 15750 10502 15802
rect 10502 15750 10554 15802
rect 10554 15750 10556 15802
rect 10180 15748 10236 15750
rect 10260 15748 10316 15750
rect 10340 15748 10396 15750
rect 10420 15748 10476 15750
rect 10500 15748 10556 15750
rect 10180 14714 10236 14716
rect 10260 14714 10316 14716
rect 10340 14714 10396 14716
rect 10420 14714 10476 14716
rect 10500 14714 10556 14716
rect 10180 14662 10182 14714
rect 10182 14662 10234 14714
rect 10234 14662 10236 14714
rect 10260 14662 10298 14714
rect 10298 14662 10310 14714
rect 10310 14662 10316 14714
rect 10340 14662 10362 14714
rect 10362 14662 10374 14714
rect 10374 14662 10396 14714
rect 10420 14662 10426 14714
rect 10426 14662 10438 14714
rect 10438 14662 10476 14714
rect 10500 14662 10502 14714
rect 10502 14662 10554 14714
rect 10554 14662 10556 14714
rect 10180 14660 10236 14662
rect 10260 14660 10316 14662
rect 10340 14660 10396 14662
rect 10420 14660 10476 14662
rect 10500 14660 10556 14662
rect 10180 13626 10236 13628
rect 10260 13626 10316 13628
rect 10340 13626 10396 13628
rect 10420 13626 10476 13628
rect 10500 13626 10556 13628
rect 10180 13574 10182 13626
rect 10182 13574 10234 13626
rect 10234 13574 10236 13626
rect 10260 13574 10298 13626
rect 10298 13574 10310 13626
rect 10310 13574 10316 13626
rect 10340 13574 10362 13626
rect 10362 13574 10374 13626
rect 10374 13574 10396 13626
rect 10420 13574 10426 13626
rect 10426 13574 10438 13626
rect 10438 13574 10476 13626
rect 10500 13574 10502 13626
rect 10502 13574 10554 13626
rect 10554 13574 10556 13626
rect 10180 13572 10236 13574
rect 10260 13572 10316 13574
rect 10340 13572 10396 13574
rect 10420 13572 10476 13574
rect 10500 13572 10556 13574
rect 10180 12538 10236 12540
rect 10260 12538 10316 12540
rect 10340 12538 10396 12540
rect 10420 12538 10476 12540
rect 10500 12538 10556 12540
rect 10180 12486 10182 12538
rect 10182 12486 10234 12538
rect 10234 12486 10236 12538
rect 10260 12486 10298 12538
rect 10298 12486 10310 12538
rect 10310 12486 10316 12538
rect 10340 12486 10362 12538
rect 10362 12486 10374 12538
rect 10374 12486 10396 12538
rect 10420 12486 10426 12538
rect 10426 12486 10438 12538
rect 10438 12486 10476 12538
rect 10500 12486 10502 12538
rect 10502 12486 10554 12538
rect 10554 12486 10556 12538
rect 10180 12484 10236 12486
rect 10260 12484 10316 12486
rect 10340 12484 10396 12486
rect 10420 12484 10476 12486
rect 10500 12484 10556 12486
rect 10180 11450 10236 11452
rect 10260 11450 10316 11452
rect 10340 11450 10396 11452
rect 10420 11450 10476 11452
rect 10500 11450 10556 11452
rect 10180 11398 10182 11450
rect 10182 11398 10234 11450
rect 10234 11398 10236 11450
rect 10260 11398 10298 11450
rect 10298 11398 10310 11450
rect 10310 11398 10316 11450
rect 10340 11398 10362 11450
rect 10362 11398 10374 11450
rect 10374 11398 10396 11450
rect 10420 11398 10426 11450
rect 10426 11398 10438 11450
rect 10438 11398 10476 11450
rect 10500 11398 10502 11450
rect 10502 11398 10554 11450
rect 10554 11398 10556 11450
rect 10180 11396 10236 11398
rect 10260 11396 10316 11398
rect 10340 11396 10396 11398
rect 10420 11396 10476 11398
rect 10500 11396 10556 11398
rect 10180 10362 10236 10364
rect 10260 10362 10316 10364
rect 10340 10362 10396 10364
rect 10420 10362 10476 10364
rect 10500 10362 10556 10364
rect 10180 10310 10182 10362
rect 10182 10310 10234 10362
rect 10234 10310 10236 10362
rect 10260 10310 10298 10362
rect 10298 10310 10310 10362
rect 10310 10310 10316 10362
rect 10340 10310 10362 10362
rect 10362 10310 10374 10362
rect 10374 10310 10396 10362
rect 10420 10310 10426 10362
rect 10426 10310 10438 10362
rect 10438 10310 10476 10362
rect 10500 10310 10502 10362
rect 10502 10310 10554 10362
rect 10554 10310 10556 10362
rect 10180 10308 10236 10310
rect 10260 10308 10316 10310
rect 10340 10308 10396 10310
rect 10420 10308 10476 10310
rect 10500 10308 10556 10310
rect 10180 9274 10236 9276
rect 10260 9274 10316 9276
rect 10340 9274 10396 9276
rect 10420 9274 10476 9276
rect 10500 9274 10556 9276
rect 10180 9222 10182 9274
rect 10182 9222 10234 9274
rect 10234 9222 10236 9274
rect 10260 9222 10298 9274
rect 10298 9222 10310 9274
rect 10310 9222 10316 9274
rect 10340 9222 10362 9274
rect 10362 9222 10374 9274
rect 10374 9222 10396 9274
rect 10420 9222 10426 9274
rect 10426 9222 10438 9274
rect 10438 9222 10476 9274
rect 10500 9222 10502 9274
rect 10502 9222 10554 9274
rect 10554 9222 10556 9274
rect 10180 9220 10236 9222
rect 10260 9220 10316 9222
rect 10340 9220 10396 9222
rect 10420 9220 10476 9222
rect 10500 9220 10556 9222
rect 9678 7420 9680 7440
rect 9680 7420 9732 7440
rect 9732 7420 9734 7440
rect 9678 7384 9734 7420
rect 4180 3834 4236 3836
rect 4260 3834 4316 3836
rect 4340 3834 4396 3836
rect 4420 3834 4476 3836
rect 4500 3834 4556 3836
rect 4180 3782 4182 3834
rect 4182 3782 4234 3834
rect 4234 3782 4236 3834
rect 4260 3782 4298 3834
rect 4298 3782 4310 3834
rect 4310 3782 4316 3834
rect 4340 3782 4362 3834
rect 4362 3782 4374 3834
rect 4374 3782 4396 3834
rect 4420 3782 4426 3834
rect 4426 3782 4438 3834
rect 4438 3782 4476 3834
rect 4500 3782 4502 3834
rect 4502 3782 4554 3834
rect 4554 3782 4556 3834
rect 4180 3780 4236 3782
rect 4260 3780 4316 3782
rect 4340 3780 4396 3782
rect 4420 3780 4476 3782
rect 4500 3780 4556 3782
rect 4920 3290 4976 3292
rect 5000 3290 5056 3292
rect 5080 3290 5136 3292
rect 5160 3290 5216 3292
rect 5240 3290 5296 3292
rect 4920 3238 4922 3290
rect 4922 3238 4974 3290
rect 4974 3238 4976 3290
rect 5000 3238 5038 3290
rect 5038 3238 5050 3290
rect 5050 3238 5056 3290
rect 5080 3238 5102 3290
rect 5102 3238 5114 3290
rect 5114 3238 5136 3290
rect 5160 3238 5166 3290
rect 5166 3238 5178 3290
rect 5178 3238 5216 3290
rect 5240 3238 5242 3290
rect 5242 3238 5294 3290
rect 5294 3238 5296 3290
rect 4920 3236 4976 3238
rect 5000 3236 5056 3238
rect 5080 3236 5136 3238
rect 5160 3236 5216 3238
rect 5240 3236 5296 3238
rect 10046 8472 10102 8528
rect 10180 8186 10236 8188
rect 10260 8186 10316 8188
rect 10340 8186 10396 8188
rect 10420 8186 10476 8188
rect 10500 8186 10556 8188
rect 10180 8134 10182 8186
rect 10182 8134 10234 8186
rect 10234 8134 10236 8186
rect 10260 8134 10298 8186
rect 10298 8134 10310 8186
rect 10310 8134 10316 8186
rect 10340 8134 10362 8186
rect 10362 8134 10374 8186
rect 10374 8134 10396 8186
rect 10420 8134 10426 8186
rect 10426 8134 10438 8186
rect 10438 8134 10476 8186
rect 10500 8134 10502 8186
rect 10502 8134 10554 8186
rect 10554 8134 10556 8186
rect 10180 8132 10236 8134
rect 10260 8132 10316 8134
rect 10340 8132 10396 8134
rect 10420 8132 10476 8134
rect 10500 8132 10556 8134
rect 9770 6704 9826 6760
rect 10180 7098 10236 7100
rect 10260 7098 10316 7100
rect 10340 7098 10396 7100
rect 10420 7098 10476 7100
rect 10500 7098 10556 7100
rect 10180 7046 10182 7098
rect 10182 7046 10234 7098
rect 10234 7046 10236 7098
rect 10260 7046 10298 7098
rect 10298 7046 10310 7098
rect 10310 7046 10316 7098
rect 10340 7046 10362 7098
rect 10362 7046 10374 7098
rect 10374 7046 10396 7098
rect 10420 7046 10426 7098
rect 10426 7046 10438 7098
rect 10438 7046 10476 7098
rect 10500 7046 10502 7098
rect 10502 7046 10554 7098
rect 10554 7046 10556 7098
rect 10180 7044 10236 7046
rect 10260 7044 10316 7046
rect 10340 7044 10396 7046
rect 10420 7044 10476 7046
rect 10500 7044 10556 7046
rect 10180 6010 10236 6012
rect 10260 6010 10316 6012
rect 10340 6010 10396 6012
rect 10420 6010 10476 6012
rect 10500 6010 10556 6012
rect 10180 5958 10182 6010
rect 10182 5958 10234 6010
rect 10234 5958 10236 6010
rect 10260 5958 10298 6010
rect 10298 5958 10310 6010
rect 10310 5958 10316 6010
rect 10340 5958 10362 6010
rect 10362 5958 10374 6010
rect 10374 5958 10396 6010
rect 10420 5958 10426 6010
rect 10426 5958 10438 6010
rect 10438 5958 10476 6010
rect 10500 5958 10502 6010
rect 10502 5958 10554 6010
rect 10554 5958 10556 6010
rect 10180 5956 10236 5958
rect 10260 5956 10316 5958
rect 10340 5956 10396 5958
rect 10420 5956 10476 5958
rect 10500 5956 10556 5958
rect 10046 4936 10102 4992
rect 10180 4922 10236 4924
rect 10260 4922 10316 4924
rect 10340 4922 10396 4924
rect 10420 4922 10476 4924
rect 10500 4922 10556 4924
rect 10180 4870 10182 4922
rect 10182 4870 10234 4922
rect 10234 4870 10236 4922
rect 10260 4870 10298 4922
rect 10298 4870 10310 4922
rect 10310 4870 10316 4922
rect 10340 4870 10362 4922
rect 10362 4870 10374 4922
rect 10374 4870 10396 4922
rect 10420 4870 10426 4922
rect 10426 4870 10438 4922
rect 10438 4870 10476 4922
rect 10500 4870 10502 4922
rect 10502 4870 10554 4922
rect 10554 4870 10556 4922
rect 10180 4868 10236 4870
rect 10260 4868 10316 4870
rect 10340 4868 10396 4870
rect 10420 4868 10476 4870
rect 10500 4868 10556 4870
rect 10920 19610 10976 19612
rect 11000 19610 11056 19612
rect 11080 19610 11136 19612
rect 11160 19610 11216 19612
rect 11240 19610 11296 19612
rect 10920 19558 10922 19610
rect 10922 19558 10974 19610
rect 10974 19558 10976 19610
rect 11000 19558 11038 19610
rect 11038 19558 11050 19610
rect 11050 19558 11056 19610
rect 11080 19558 11102 19610
rect 11102 19558 11114 19610
rect 11114 19558 11136 19610
rect 11160 19558 11166 19610
rect 11166 19558 11178 19610
rect 11178 19558 11216 19610
rect 11240 19558 11242 19610
rect 11242 19558 11294 19610
rect 11294 19558 11296 19610
rect 10920 19556 10976 19558
rect 11000 19556 11056 19558
rect 11080 19556 11136 19558
rect 11160 19556 11216 19558
rect 11240 19556 11296 19558
rect 12162 20712 12218 20768
rect 10920 18522 10976 18524
rect 11000 18522 11056 18524
rect 11080 18522 11136 18524
rect 11160 18522 11216 18524
rect 11240 18522 11296 18524
rect 10920 18470 10922 18522
rect 10922 18470 10974 18522
rect 10974 18470 10976 18522
rect 11000 18470 11038 18522
rect 11038 18470 11050 18522
rect 11050 18470 11056 18522
rect 11080 18470 11102 18522
rect 11102 18470 11114 18522
rect 11114 18470 11136 18522
rect 11160 18470 11166 18522
rect 11166 18470 11178 18522
rect 11178 18470 11216 18522
rect 11240 18470 11242 18522
rect 11242 18470 11294 18522
rect 11294 18470 11296 18522
rect 10920 18468 10976 18470
rect 11000 18468 11056 18470
rect 11080 18468 11136 18470
rect 11160 18468 11216 18470
rect 11240 18468 11296 18470
rect 10920 17434 10976 17436
rect 11000 17434 11056 17436
rect 11080 17434 11136 17436
rect 11160 17434 11216 17436
rect 11240 17434 11296 17436
rect 10920 17382 10922 17434
rect 10922 17382 10974 17434
rect 10974 17382 10976 17434
rect 11000 17382 11038 17434
rect 11038 17382 11050 17434
rect 11050 17382 11056 17434
rect 11080 17382 11102 17434
rect 11102 17382 11114 17434
rect 11114 17382 11136 17434
rect 11160 17382 11166 17434
rect 11166 17382 11178 17434
rect 11178 17382 11216 17434
rect 11240 17382 11242 17434
rect 11242 17382 11294 17434
rect 11294 17382 11296 17434
rect 10920 17380 10976 17382
rect 11000 17380 11056 17382
rect 11080 17380 11136 17382
rect 11160 17380 11216 17382
rect 11240 17380 11296 17382
rect 10920 16346 10976 16348
rect 11000 16346 11056 16348
rect 11080 16346 11136 16348
rect 11160 16346 11216 16348
rect 11240 16346 11296 16348
rect 10920 16294 10922 16346
rect 10922 16294 10974 16346
rect 10974 16294 10976 16346
rect 11000 16294 11038 16346
rect 11038 16294 11050 16346
rect 11050 16294 11056 16346
rect 11080 16294 11102 16346
rect 11102 16294 11114 16346
rect 11114 16294 11136 16346
rect 11160 16294 11166 16346
rect 11166 16294 11178 16346
rect 11178 16294 11216 16346
rect 11240 16294 11242 16346
rect 11242 16294 11294 16346
rect 11294 16294 11296 16346
rect 10920 16292 10976 16294
rect 11000 16292 11056 16294
rect 11080 16292 11136 16294
rect 11160 16292 11216 16294
rect 11240 16292 11296 16294
rect 10920 15258 10976 15260
rect 11000 15258 11056 15260
rect 11080 15258 11136 15260
rect 11160 15258 11216 15260
rect 11240 15258 11296 15260
rect 10920 15206 10922 15258
rect 10922 15206 10974 15258
rect 10974 15206 10976 15258
rect 11000 15206 11038 15258
rect 11038 15206 11050 15258
rect 11050 15206 11056 15258
rect 11080 15206 11102 15258
rect 11102 15206 11114 15258
rect 11114 15206 11136 15258
rect 11160 15206 11166 15258
rect 11166 15206 11178 15258
rect 11178 15206 11216 15258
rect 11240 15206 11242 15258
rect 11242 15206 11294 15258
rect 11294 15206 11296 15258
rect 10920 15204 10976 15206
rect 11000 15204 11056 15206
rect 11080 15204 11136 15206
rect 11160 15204 11216 15206
rect 11240 15204 11296 15206
rect 10920 14170 10976 14172
rect 11000 14170 11056 14172
rect 11080 14170 11136 14172
rect 11160 14170 11216 14172
rect 11240 14170 11296 14172
rect 10920 14118 10922 14170
rect 10922 14118 10974 14170
rect 10974 14118 10976 14170
rect 11000 14118 11038 14170
rect 11038 14118 11050 14170
rect 11050 14118 11056 14170
rect 11080 14118 11102 14170
rect 11102 14118 11114 14170
rect 11114 14118 11136 14170
rect 11160 14118 11166 14170
rect 11166 14118 11178 14170
rect 11178 14118 11216 14170
rect 11240 14118 11242 14170
rect 11242 14118 11294 14170
rect 11294 14118 11296 14170
rect 10920 14116 10976 14118
rect 11000 14116 11056 14118
rect 11080 14116 11136 14118
rect 11160 14116 11216 14118
rect 11240 14116 11296 14118
rect 10920 13082 10976 13084
rect 11000 13082 11056 13084
rect 11080 13082 11136 13084
rect 11160 13082 11216 13084
rect 11240 13082 11296 13084
rect 10920 13030 10922 13082
rect 10922 13030 10974 13082
rect 10974 13030 10976 13082
rect 11000 13030 11038 13082
rect 11038 13030 11050 13082
rect 11050 13030 11056 13082
rect 11080 13030 11102 13082
rect 11102 13030 11114 13082
rect 11114 13030 11136 13082
rect 11160 13030 11166 13082
rect 11166 13030 11178 13082
rect 11178 13030 11216 13082
rect 11240 13030 11242 13082
rect 11242 13030 11294 13082
rect 11294 13030 11296 13082
rect 10920 13028 10976 13030
rect 11000 13028 11056 13030
rect 11080 13028 11136 13030
rect 11160 13028 11216 13030
rect 11240 13028 11296 13030
rect 10920 11994 10976 11996
rect 11000 11994 11056 11996
rect 11080 11994 11136 11996
rect 11160 11994 11216 11996
rect 11240 11994 11296 11996
rect 10920 11942 10922 11994
rect 10922 11942 10974 11994
rect 10974 11942 10976 11994
rect 11000 11942 11038 11994
rect 11038 11942 11050 11994
rect 11050 11942 11056 11994
rect 11080 11942 11102 11994
rect 11102 11942 11114 11994
rect 11114 11942 11136 11994
rect 11160 11942 11166 11994
rect 11166 11942 11178 11994
rect 11178 11942 11216 11994
rect 11240 11942 11242 11994
rect 11242 11942 11294 11994
rect 11294 11942 11296 11994
rect 10920 11940 10976 11942
rect 11000 11940 11056 11942
rect 11080 11940 11136 11942
rect 11160 11940 11216 11942
rect 11240 11940 11296 11942
rect 10920 10906 10976 10908
rect 11000 10906 11056 10908
rect 11080 10906 11136 10908
rect 11160 10906 11216 10908
rect 11240 10906 11296 10908
rect 10920 10854 10922 10906
rect 10922 10854 10974 10906
rect 10974 10854 10976 10906
rect 11000 10854 11038 10906
rect 11038 10854 11050 10906
rect 11050 10854 11056 10906
rect 11080 10854 11102 10906
rect 11102 10854 11114 10906
rect 11114 10854 11136 10906
rect 11160 10854 11166 10906
rect 11166 10854 11178 10906
rect 11178 10854 11216 10906
rect 11240 10854 11242 10906
rect 11242 10854 11294 10906
rect 11294 10854 11296 10906
rect 10920 10852 10976 10854
rect 11000 10852 11056 10854
rect 11080 10852 11136 10854
rect 11160 10852 11216 10854
rect 11240 10852 11296 10854
rect 10920 9818 10976 9820
rect 11000 9818 11056 9820
rect 11080 9818 11136 9820
rect 11160 9818 11216 9820
rect 11240 9818 11296 9820
rect 10920 9766 10922 9818
rect 10922 9766 10974 9818
rect 10974 9766 10976 9818
rect 11000 9766 11038 9818
rect 11038 9766 11050 9818
rect 11050 9766 11056 9818
rect 11080 9766 11102 9818
rect 11102 9766 11114 9818
rect 11114 9766 11136 9818
rect 11160 9766 11166 9818
rect 11166 9766 11178 9818
rect 11178 9766 11216 9818
rect 11240 9766 11242 9818
rect 11242 9766 11294 9818
rect 11294 9766 11296 9818
rect 10920 9764 10976 9766
rect 11000 9764 11056 9766
rect 11080 9764 11136 9766
rect 11160 9764 11216 9766
rect 11240 9764 11296 9766
rect 10782 8880 10838 8936
rect 10920 8730 10976 8732
rect 11000 8730 11056 8732
rect 11080 8730 11136 8732
rect 11160 8730 11216 8732
rect 11240 8730 11296 8732
rect 10920 8678 10922 8730
rect 10922 8678 10974 8730
rect 10974 8678 10976 8730
rect 11000 8678 11038 8730
rect 11038 8678 11050 8730
rect 11050 8678 11056 8730
rect 11080 8678 11102 8730
rect 11102 8678 11114 8730
rect 11114 8678 11136 8730
rect 11160 8678 11166 8730
rect 11166 8678 11178 8730
rect 11178 8678 11216 8730
rect 11240 8678 11242 8730
rect 11242 8678 11294 8730
rect 11294 8678 11296 8730
rect 10920 8676 10976 8678
rect 11000 8676 11056 8678
rect 11080 8676 11136 8678
rect 11160 8676 11216 8678
rect 11240 8676 11296 8678
rect 22180 32122 22236 32124
rect 22260 32122 22316 32124
rect 22340 32122 22396 32124
rect 22420 32122 22476 32124
rect 22500 32122 22556 32124
rect 22180 32070 22182 32122
rect 22182 32070 22234 32122
rect 22234 32070 22236 32122
rect 22260 32070 22298 32122
rect 22298 32070 22310 32122
rect 22310 32070 22316 32122
rect 22340 32070 22362 32122
rect 22362 32070 22374 32122
rect 22374 32070 22396 32122
rect 22420 32070 22426 32122
rect 22426 32070 22438 32122
rect 22438 32070 22476 32122
rect 22500 32070 22502 32122
rect 22502 32070 22554 32122
rect 22554 32070 22556 32122
rect 22180 32068 22236 32070
rect 22260 32068 22316 32070
rect 22340 32068 22396 32070
rect 22420 32068 22476 32070
rect 22500 32068 22556 32070
rect 16920 31578 16976 31580
rect 17000 31578 17056 31580
rect 17080 31578 17136 31580
rect 17160 31578 17216 31580
rect 17240 31578 17296 31580
rect 16920 31526 16922 31578
rect 16922 31526 16974 31578
rect 16974 31526 16976 31578
rect 17000 31526 17038 31578
rect 17038 31526 17050 31578
rect 17050 31526 17056 31578
rect 17080 31526 17102 31578
rect 17102 31526 17114 31578
rect 17114 31526 17136 31578
rect 17160 31526 17166 31578
rect 17166 31526 17178 31578
rect 17178 31526 17216 31578
rect 17240 31526 17242 31578
rect 17242 31526 17294 31578
rect 17294 31526 17296 31578
rect 16920 31524 16976 31526
rect 17000 31524 17056 31526
rect 17080 31524 17136 31526
rect 17160 31524 17216 31526
rect 17240 31524 17296 31526
rect 16180 31034 16236 31036
rect 16260 31034 16316 31036
rect 16340 31034 16396 31036
rect 16420 31034 16476 31036
rect 16500 31034 16556 31036
rect 16180 30982 16182 31034
rect 16182 30982 16234 31034
rect 16234 30982 16236 31034
rect 16260 30982 16298 31034
rect 16298 30982 16310 31034
rect 16310 30982 16316 31034
rect 16340 30982 16362 31034
rect 16362 30982 16374 31034
rect 16374 30982 16396 31034
rect 16420 30982 16426 31034
rect 16426 30982 16438 31034
rect 16438 30982 16476 31034
rect 16500 30982 16502 31034
rect 16502 30982 16554 31034
rect 16554 30982 16556 31034
rect 16180 30980 16236 30982
rect 16260 30980 16316 30982
rect 16340 30980 16396 30982
rect 16420 30980 16476 30982
rect 16500 30980 16556 30982
rect 14002 29008 14058 29064
rect 14094 23432 14150 23488
rect 16180 29946 16236 29948
rect 16260 29946 16316 29948
rect 16340 29946 16396 29948
rect 16420 29946 16476 29948
rect 16500 29946 16556 29948
rect 16180 29894 16182 29946
rect 16182 29894 16234 29946
rect 16234 29894 16236 29946
rect 16260 29894 16298 29946
rect 16298 29894 16310 29946
rect 16310 29894 16316 29946
rect 16340 29894 16362 29946
rect 16362 29894 16374 29946
rect 16374 29894 16396 29946
rect 16420 29894 16426 29946
rect 16426 29894 16438 29946
rect 16438 29894 16476 29946
rect 16500 29894 16502 29946
rect 16502 29894 16554 29946
rect 16554 29894 16556 29946
rect 16180 29892 16236 29894
rect 16260 29892 16316 29894
rect 16340 29892 16396 29894
rect 16420 29892 16476 29894
rect 16500 29892 16556 29894
rect 10920 7642 10976 7644
rect 11000 7642 11056 7644
rect 11080 7642 11136 7644
rect 11160 7642 11216 7644
rect 11240 7642 11296 7644
rect 10920 7590 10922 7642
rect 10922 7590 10974 7642
rect 10974 7590 10976 7642
rect 11000 7590 11038 7642
rect 11038 7590 11050 7642
rect 11050 7590 11056 7642
rect 11080 7590 11102 7642
rect 11102 7590 11114 7642
rect 11114 7590 11136 7642
rect 11160 7590 11166 7642
rect 11166 7590 11178 7642
rect 11178 7590 11216 7642
rect 11240 7590 11242 7642
rect 11242 7590 11294 7642
rect 11294 7590 11296 7642
rect 10920 7588 10976 7590
rect 11000 7588 11056 7590
rect 11080 7588 11136 7590
rect 11160 7588 11216 7590
rect 11240 7588 11296 7590
rect 10920 6554 10976 6556
rect 11000 6554 11056 6556
rect 11080 6554 11136 6556
rect 11160 6554 11216 6556
rect 11240 6554 11296 6556
rect 10920 6502 10922 6554
rect 10922 6502 10974 6554
rect 10974 6502 10976 6554
rect 11000 6502 11038 6554
rect 11038 6502 11050 6554
rect 11050 6502 11056 6554
rect 11080 6502 11102 6554
rect 11102 6502 11114 6554
rect 11114 6502 11136 6554
rect 11160 6502 11166 6554
rect 11166 6502 11178 6554
rect 11178 6502 11216 6554
rect 11240 6502 11242 6554
rect 11242 6502 11294 6554
rect 11294 6502 11296 6554
rect 10920 6500 10976 6502
rect 11000 6500 11056 6502
rect 11080 6500 11136 6502
rect 11160 6500 11216 6502
rect 11240 6500 11296 6502
rect 12990 11328 13046 11384
rect 14370 19388 14372 19408
rect 14372 19388 14424 19408
rect 14424 19388 14426 19408
rect 14370 19352 14426 19388
rect 16920 30490 16976 30492
rect 17000 30490 17056 30492
rect 17080 30490 17136 30492
rect 17160 30490 17216 30492
rect 17240 30490 17296 30492
rect 16920 30438 16922 30490
rect 16922 30438 16974 30490
rect 16974 30438 16976 30490
rect 17000 30438 17038 30490
rect 17038 30438 17050 30490
rect 17050 30438 17056 30490
rect 17080 30438 17102 30490
rect 17102 30438 17114 30490
rect 17114 30438 17136 30490
rect 17160 30438 17166 30490
rect 17166 30438 17178 30490
rect 17178 30438 17216 30490
rect 17240 30438 17242 30490
rect 17242 30438 17294 30490
rect 17294 30438 17296 30490
rect 16920 30436 16976 30438
rect 17000 30436 17056 30438
rect 17080 30436 17136 30438
rect 17160 30436 17216 30438
rect 17240 30436 17296 30438
rect 16180 28858 16236 28860
rect 16260 28858 16316 28860
rect 16340 28858 16396 28860
rect 16420 28858 16476 28860
rect 16500 28858 16556 28860
rect 16180 28806 16182 28858
rect 16182 28806 16234 28858
rect 16234 28806 16236 28858
rect 16260 28806 16298 28858
rect 16298 28806 16310 28858
rect 16310 28806 16316 28858
rect 16340 28806 16362 28858
rect 16362 28806 16374 28858
rect 16374 28806 16396 28858
rect 16420 28806 16426 28858
rect 16426 28806 16438 28858
rect 16438 28806 16476 28858
rect 16500 28806 16502 28858
rect 16502 28806 16554 28858
rect 16554 28806 16556 28858
rect 16180 28804 16236 28806
rect 16260 28804 16316 28806
rect 16340 28804 16396 28806
rect 16420 28804 16476 28806
rect 16500 28804 16556 28806
rect 16920 29402 16976 29404
rect 17000 29402 17056 29404
rect 17080 29402 17136 29404
rect 17160 29402 17216 29404
rect 17240 29402 17296 29404
rect 16920 29350 16922 29402
rect 16922 29350 16974 29402
rect 16974 29350 16976 29402
rect 17000 29350 17038 29402
rect 17038 29350 17050 29402
rect 17050 29350 17056 29402
rect 17080 29350 17102 29402
rect 17102 29350 17114 29402
rect 17114 29350 17136 29402
rect 17160 29350 17166 29402
rect 17166 29350 17178 29402
rect 17178 29350 17216 29402
rect 17240 29350 17242 29402
rect 17242 29350 17294 29402
rect 17294 29350 17296 29402
rect 16920 29348 16976 29350
rect 17000 29348 17056 29350
rect 17080 29348 17136 29350
rect 17160 29348 17216 29350
rect 17240 29348 17296 29350
rect 16920 28314 16976 28316
rect 17000 28314 17056 28316
rect 17080 28314 17136 28316
rect 17160 28314 17216 28316
rect 17240 28314 17296 28316
rect 16920 28262 16922 28314
rect 16922 28262 16974 28314
rect 16974 28262 16976 28314
rect 17000 28262 17038 28314
rect 17038 28262 17050 28314
rect 17050 28262 17056 28314
rect 17080 28262 17102 28314
rect 17102 28262 17114 28314
rect 17114 28262 17136 28314
rect 17160 28262 17166 28314
rect 17166 28262 17178 28314
rect 17178 28262 17216 28314
rect 17240 28262 17242 28314
rect 17242 28262 17294 28314
rect 17294 28262 17296 28314
rect 16920 28260 16976 28262
rect 17000 28260 17056 28262
rect 17080 28260 17136 28262
rect 17160 28260 17216 28262
rect 17240 28260 17296 28262
rect 16180 27770 16236 27772
rect 16260 27770 16316 27772
rect 16340 27770 16396 27772
rect 16420 27770 16476 27772
rect 16500 27770 16556 27772
rect 16180 27718 16182 27770
rect 16182 27718 16234 27770
rect 16234 27718 16236 27770
rect 16260 27718 16298 27770
rect 16298 27718 16310 27770
rect 16310 27718 16316 27770
rect 16340 27718 16362 27770
rect 16362 27718 16374 27770
rect 16374 27718 16396 27770
rect 16420 27718 16426 27770
rect 16426 27718 16438 27770
rect 16438 27718 16476 27770
rect 16500 27718 16502 27770
rect 16502 27718 16554 27770
rect 16554 27718 16556 27770
rect 16180 27716 16236 27718
rect 16260 27716 16316 27718
rect 16340 27716 16396 27718
rect 16420 27716 16476 27718
rect 16500 27716 16556 27718
rect 15934 27376 15990 27432
rect 16118 26832 16174 26888
rect 16180 26682 16236 26684
rect 16260 26682 16316 26684
rect 16340 26682 16396 26684
rect 16420 26682 16476 26684
rect 16500 26682 16556 26684
rect 16180 26630 16182 26682
rect 16182 26630 16234 26682
rect 16234 26630 16236 26682
rect 16260 26630 16298 26682
rect 16298 26630 16310 26682
rect 16310 26630 16316 26682
rect 16340 26630 16362 26682
rect 16362 26630 16374 26682
rect 16374 26630 16396 26682
rect 16420 26630 16426 26682
rect 16426 26630 16438 26682
rect 16438 26630 16476 26682
rect 16500 26630 16502 26682
rect 16502 26630 16554 26682
rect 16554 26630 16556 26682
rect 16180 26628 16236 26630
rect 16260 26628 16316 26630
rect 16340 26628 16396 26630
rect 16420 26628 16476 26630
rect 16500 26628 16556 26630
rect 16920 27226 16976 27228
rect 17000 27226 17056 27228
rect 17080 27226 17136 27228
rect 17160 27226 17216 27228
rect 17240 27226 17296 27228
rect 16920 27174 16922 27226
rect 16922 27174 16974 27226
rect 16974 27174 16976 27226
rect 17000 27174 17038 27226
rect 17038 27174 17050 27226
rect 17050 27174 17056 27226
rect 17080 27174 17102 27226
rect 17102 27174 17114 27226
rect 17114 27174 17136 27226
rect 17160 27174 17166 27226
rect 17166 27174 17178 27226
rect 17178 27174 17216 27226
rect 17240 27174 17242 27226
rect 17242 27174 17294 27226
rect 17294 27174 17296 27226
rect 16920 27172 16976 27174
rect 17000 27172 17056 27174
rect 17080 27172 17136 27174
rect 17160 27172 17216 27174
rect 17240 27172 17296 27174
rect 16854 26696 16910 26752
rect 17130 26832 17186 26888
rect 17774 27376 17830 27432
rect 16920 26138 16976 26140
rect 17000 26138 17056 26140
rect 17080 26138 17136 26140
rect 17160 26138 17216 26140
rect 17240 26138 17296 26140
rect 16920 26086 16922 26138
rect 16922 26086 16974 26138
rect 16974 26086 16976 26138
rect 17000 26086 17038 26138
rect 17038 26086 17050 26138
rect 17050 26086 17056 26138
rect 17080 26086 17102 26138
rect 17102 26086 17114 26138
rect 17114 26086 17136 26138
rect 17160 26086 17166 26138
rect 17166 26086 17178 26138
rect 17178 26086 17216 26138
rect 17240 26086 17242 26138
rect 17242 26086 17294 26138
rect 17294 26086 17296 26138
rect 16920 26084 16976 26086
rect 17000 26084 17056 26086
rect 17080 26084 17136 26086
rect 17160 26084 17216 26086
rect 17240 26084 17296 26086
rect 16180 25594 16236 25596
rect 16260 25594 16316 25596
rect 16340 25594 16396 25596
rect 16420 25594 16476 25596
rect 16500 25594 16556 25596
rect 16180 25542 16182 25594
rect 16182 25542 16234 25594
rect 16234 25542 16236 25594
rect 16260 25542 16298 25594
rect 16298 25542 16310 25594
rect 16310 25542 16316 25594
rect 16340 25542 16362 25594
rect 16362 25542 16374 25594
rect 16374 25542 16396 25594
rect 16420 25542 16426 25594
rect 16426 25542 16438 25594
rect 16438 25542 16476 25594
rect 16500 25542 16502 25594
rect 16502 25542 16554 25594
rect 16554 25542 16556 25594
rect 16180 25540 16236 25542
rect 16260 25540 16316 25542
rect 16340 25540 16396 25542
rect 16420 25540 16476 25542
rect 16500 25540 16556 25542
rect 16920 25050 16976 25052
rect 17000 25050 17056 25052
rect 17080 25050 17136 25052
rect 17160 25050 17216 25052
rect 17240 25050 17296 25052
rect 16920 24998 16922 25050
rect 16922 24998 16974 25050
rect 16974 24998 16976 25050
rect 17000 24998 17038 25050
rect 17038 24998 17050 25050
rect 17050 24998 17056 25050
rect 17080 24998 17102 25050
rect 17102 24998 17114 25050
rect 17114 24998 17136 25050
rect 17160 24998 17166 25050
rect 17166 24998 17178 25050
rect 17178 24998 17216 25050
rect 17240 24998 17242 25050
rect 17242 24998 17294 25050
rect 17294 24998 17296 25050
rect 16920 24996 16976 24998
rect 17000 24996 17056 24998
rect 17080 24996 17136 24998
rect 17160 24996 17216 24998
rect 17240 24996 17296 24998
rect 18050 26832 18106 26888
rect 18326 26696 18382 26752
rect 16180 24506 16236 24508
rect 16260 24506 16316 24508
rect 16340 24506 16396 24508
rect 16420 24506 16476 24508
rect 16500 24506 16556 24508
rect 16180 24454 16182 24506
rect 16182 24454 16234 24506
rect 16234 24454 16236 24506
rect 16260 24454 16298 24506
rect 16298 24454 16310 24506
rect 16310 24454 16316 24506
rect 16340 24454 16362 24506
rect 16362 24454 16374 24506
rect 16374 24454 16396 24506
rect 16420 24454 16426 24506
rect 16426 24454 16438 24506
rect 16438 24454 16476 24506
rect 16500 24454 16502 24506
rect 16502 24454 16554 24506
rect 16554 24454 16556 24506
rect 16180 24452 16236 24454
rect 16260 24452 16316 24454
rect 16340 24452 16396 24454
rect 16420 24452 16476 24454
rect 16500 24452 16556 24454
rect 16920 23962 16976 23964
rect 17000 23962 17056 23964
rect 17080 23962 17136 23964
rect 17160 23962 17216 23964
rect 17240 23962 17296 23964
rect 16920 23910 16922 23962
rect 16922 23910 16974 23962
rect 16974 23910 16976 23962
rect 17000 23910 17038 23962
rect 17038 23910 17050 23962
rect 17050 23910 17056 23962
rect 17080 23910 17102 23962
rect 17102 23910 17114 23962
rect 17114 23910 17136 23962
rect 17160 23910 17166 23962
rect 17166 23910 17178 23962
rect 17178 23910 17216 23962
rect 17240 23910 17242 23962
rect 17242 23910 17294 23962
rect 17294 23910 17296 23962
rect 16920 23908 16976 23910
rect 17000 23908 17056 23910
rect 17080 23908 17136 23910
rect 17160 23908 17216 23910
rect 17240 23908 17296 23910
rect 16180 23418 16236 23420
rect 16260 23418 16316 23420
rect 16340 23418 16396 23420
rect 16420 23418 16476 23420
rect 16500 23418 16556 23420
rect 16180 23366 16182 23418
rect 16182 23366 16234 23418
rect 16234 23366 16236 23418
rect 16260 23366 16298 23418
rect 16298 23366 16310 23418
rect 16310 23366 16316 23418
rect 16340 23366 16362 23418
rect 16362 23366 16374 23418
rect 16374 23366 16396 23418
rect 16420 23366 16426 23418
rect 16426 23366 16438 23418
rect 16438 23366 16476 23418
rect 16500 23366 16502 23418
rect 16502 23366 16554 23418
rect 16554 23366 16556 23418
rect 16180 23364 16236 23366
rect 16260 23364 16316 23366
rect 16340 23364 16396 23366
rect 16420 23364 16476 23366
rect 16500 23364 16556 23366
rect 16920 22874 16976 22876
rect 17000 22874 17056 22876
rect 17080 22874 17136 22876
rect 17160 22874 17216 22876
rect 17240 22874 17296 22876
rect 16920 22822 16922 22874
rect 16922 22822 16974 22874
rect 16974 22822 16976 22874
rect 17000 22822 17038 22874
rect 17038 22822 17050 22874
rect 17050 22822 17056 22874
rect 17080 22822 17102 22874
rect 17102 22822 17114 22874
rect 17114 22822 17136 22874
rect 17160 22822 17166 22874
rect 17166 22822 17178 22874
rect 17178 22822 17216 22874
rect 17240 22822 17242 22874
rect 17242 22822 17294 22874
rect 17294 22822 17296 22874
rect 16920 22820 16976 22822
rect 17000 22820 17056 22822
rect 17080 22820 17136 22822
rect 17160 22820 17216 22822
rect 17240 22820 17296 22822
rect 16180 22330 16236 22332
rect 16260 22330 16316 22332
rect 16340 22330 16396 22332
rect 16420 22330 16476 22332
rect 16500 22330 16556 22332
rect 16180 22278 16182 22330
rect 16182 22278 16234 22330
rect 16234 22278 16236 22330
rect 16260 22278 16298 22330
rect 16298 22278 16310 22330
rect 16310 22278 16316 22330
rect 16340 22278 16362 22330
rect 16362 22278 16374 22330
rect 16374 22278 16396 22330
rect 16420 22278 16426 22330
rect 16426 22278 16438 22330
rect 16438 22278 16476 22330
rect 16500 22278 16502 22330
rect 16502 22278 16554 22330
rect 16554 22278 16556 22330
rect 16180 22276 16236 22278
rect 16260 22276 16316 22278
rect 16340 22276 16396 22278
rect 16420 22276 16476 22278
rect 16500 22276 16556 22278
rect 16920 21786 16976 21788
rect 17000 21786 17056 21788
rect 17080 21786 17136 21788
rect 17160 21786 17216 21788
rect 17240 21786 17296 21788
rect 16920 21734 16922 21786
rect 16922 21734 16974 21786
rect 16974 21734 16976 21786
rect 17000 21734 17038 21786
rect 17038 21734 17050 21786
rect 17050 21734 17056 21786
rect 17080 21734 17102 21786
rect 17102 21734 17114 21786
rect 17114 21734 17136 21786
rect 17160 21734 17166 21786
rect 17166 21734 17178 21786
rect 17178 21734 17216 21786
rect 17240 21734 17242 21786
rect 17242 21734 17294 21786
rect 17294 21734 17296 21786
rect 16920 21732 16976 21734
rect 17000 21732 17056 21734
rect 17080 21732 17136 21734
rect 17160 21732 17216 21734
rect 17240 21732 17296 21734
rect 22920 31578 22976 31580
rect 23000 31578 23056 31580
rect 23080 31578 23136 31580
rect 23160 31578 23216 31580
rect 23240 31578 23296 31580
rect 22920 31526 22922 31578
rect 22922 31526 22974 31578
rect 22974 31526 22976 31578
rect 23000 31526 23038 31578
rect 23038 31526 23050 31578
rect 23050 31526 23056 31578
rect 23080 31526 23102 31578
rect 23102 31526 23114 31578
rect 23114 31526 23136 31578
rect 23160 31526 23166 31578
rect 23166 31526 23178 31578
rect 23178 31526 23216 31578
rect 23240 31526 23242 31578
rect 23242 31526 23294 31578
rect 23294 31526 23296 31578
rect 22920 31524 22976 31526
rect 23000 31524 23056 31526
rect 23080 31524 23136 31526
rect 23160 31524 23216 31526
rect 23240 31524 23296 31526
rect 28180 32122 28236 32124
rect 28260 32122 28316 32124
rect 28340 32122 28396 32124
rect 28420 32122 28476 32124
rect 28500 32122 28556 32124
rect 28180 32070 28182 32122
rect 28182 32070 28234 32122
rect 28234 32070 28236 32122
rect 28260 32070 28298 32122
rect 28298 32070 28310 32122
rect 28310 32070 28316 32122
rect 28340 32070 28362 32122
rect 28362 32070 28374 32122
rect 28374 32070 28396 32122
rect 28420 32070 28426 32122
rect 28426 32070 28438 32122
rect 28438 32070 28476 32122
rect 28500 32070 28502 32122
rect 28502 32070 28554 32122
rect 28554 32070 28556 32122
rect 28180 32068 28236 32070
rect 28260 32068 28316 32070
rect 28340 32068 28396 32070
rect 28420 32068 28476 32070
rect 28500 32068 28556 32070
rect 28920 31578 28976 31580
rect 29000 31578 29056 31580
rect 29080 31578 29136 31580
rect 29160 31578 29216 31580
rect 29240 31578 29296 31580
rect 28920 31526 28922 31578
rect 28922 31526 28974 31578
rect 28974 31526 28976 31578
rect 29000 31526 29038 31578
rect 29038 31526 29050 31578
rect 29050 31526 29056 31578
rect 29080 31526 29102 31578
rect 29102 31526 29114 31578
rect 29114 31526 29136 31578
rect 29160 31526 29166 31578
rect 29166 31526 29178 31578
rect 29178 31526 29216 31578
rect 29240 31526 29242 31578
rect 29242 31526 29294 31578
rect 29294 31526 29296 31578
rect 28920 31524 28976 31526
rect 29000 31524 29056 31526
rect 29080 31524 29136 31526
rect 29160 31524 29216 31526
rect 29240 31524 29296 31526
rect 22180 31034 22236 31036
rect 22260 31034 22316 31036
rect 22340 31034 22396 31036
rect 22420 31034 22476 31036
rect 22500 31034 22556 31036
rect 22180 30982 22182 31034
rect 22182 30982 22234 31034
rect 22234 30982 22236 31034
rect 22260 30982 22298 31034
rect 22298 30982 22310 31034
rect 22310 30982 22316 31034
rect 22340 30982 22362 31034
rect 22362 30982 22374 31034
rect 22374 30982 22396 31034
rect 22420 30982 22426 31034
rect 22426 30982 22438 31034
rect 22438 30982 22476 31034
rect 22500 30982 22502 31034
rect 22502 30982 22554 31034
rect 22554 30982 22556 31034
rect 22180 30980 22236 30982
rect 22260 30980 22316 30982
rect 22340 30980 22396 30982
rect 22420 30980 22476 30982
rect 22500 30980 22556 30982
rect 28180 31034 28236 31036
rect 28260 31034 28316 31036
rect 28340 31034 28396 31036
rect 28420 31034 28476 31036
rect 28500 31034 28556 31036
rect 28180 30982 28182 31034
rect 28182 30982 28234 31034
rect 28234 30982 28236 31034
rect 28260 30982 28298 31034
rect 28298 30982 28310 31034
rect 28310 30982 28316 31034
rect 28340 30982 28362 31034
rect 28362 30982 28374 31034
rect 28374 30982 28396 31034
rect 28420 30982 28426 31034
rect 28426 30982 28438 31034
rect 28438 30982 28476 31034
rect 28500 30982 28502 31034
rect 28502 30982 28554 31034
rect 28554 30982 28556 31034
rect 28180 30980 28236 30982
rect 28260 30980 28316 30982
rect 28340 30980 28396 30982
rect 28420 30980 28476 30982
rect 28500 30980 28556 30982
rect 22920 30490 22976 30492
rect 23000 30490 23056 30492
rect 23080 30490 23136 30492
rect 23160 30490 23216 30492
rect 23240 30490 23296 30492
rect 22920 30438 22922 30490
rect 22922 30438 22974 30490
rect 22974 30438 22976 30490
rect 23000 30438 23038 30490
rect 23038 30438 23050 30490
rect 23050 30438 23056 30490
rect 23080 30438 23102 30490
rect 23102 30438 23114 30490
rect 23114 30438 23136 30490
rect 23160 30438 23166 30490
rect 23166 30438 23178 30490
rect 23178 30438 23216 30490
rect 23240 30438 23242 30490
rect 23242 30438 23294 30490
rect 23294 30438 23296 30490
rect 22920 30436 22976 30438
rect 23000 30436 23056 30438
rect 23080 30436 23136 30438
rect 23160 30436 23216 30438
rect 23240 30436 23296 30438
rect 28920 30490 28976 30492
rect 29000 30490 29056 30492
rect 29080 30490 29136 30492
rect 29160 30490 29216 30492
rect 29240 30490 29296 30492
rect 28920 30438 28922 30490
rect 28922 30438 28974 30490
rect 28974 30438 28976 30490
rect 29000 30438 29038 30490
rect 29038 30438 29050 30490
rect 29050 30438 29056 30490
rect 29080 30438 29102 30490
rect 29102 30438 29114 30490
rect 29114 30438 29136 30490
rect 29160 30438 29166 30490
rect 29166 30438 29178 30490
rect 29178 30438 29216 30490
rect 29240 30438 29242 30490
rect 29242 30438 29294 30490
rect 29294 30438 29296 30490
rect 28920 30436 28976 30438
rect 29000 30436 29056 30438
rect 29080 30436 29136 30438
rect 29160 30436 29216 30438
rect 29240 30436 29296 30438
rect 22180 29946 22236 29948
rect 22260 29946 22316 29948
rect 22340 29946 22396 29948
rect 22420 29946 22476 29948
rect 22500 29946 22556 29948
rect 22180 29894 22182 29946
rect 22182 29894 22234 29946
rect 22234 29894 22236 29946
rect 22260 29894 22298 29946
rect 22298 29894 22310 29946
rect 22310 29894 22316 29946
rect 22340 29894 22362 29946
rect 22362 29894 22374 29946
rect 22374 29894 22396 29946
rect 22420 29894 22426 29946
rect 22426 29894 22438 29946
rect 22438 29894 22476 29946
rect 22500 29894 22502 29946
rect 22502 29894 22554 29946
rect 22554 29894 22556 29946
rect 22180 29892 22236 29894
rect 22260 29892 22316 29894
rect 22340 29892 22396 29894
rect 22420 29892 22476 29894
rect 22500 29892 22556 29894
rect 28180 29946 28236 29948
rect 28260 29946 28316 29948
rect 28340 29946 28396 29948
rect 28420 29946 28476 29948
rect 28500 29946 28556 29948
rect 28180 29894 28182 29946
rect 28182 29894 28234 29946
rect 28234 29894 28236 29946
rect 28260 29894 28298 29946
rect 28298 29894 28310 29946
rect 28310 29894 28316 29946
rect 28340 29894 28362 29946
rect 28362 29894 28374 29946
rect 28374 29894 28396 29946
rect 28420 29894 28426 29946
rect 28426 29894 28438 29946
rect 28438 29894 28476 29946
rect 28500 29894 28502 29946
rect 28502 29894 28554 29946
rect 28554 29894 28556 29946
rect 28180 29892 28236 29894
rect 28260 29892 28316 29894
rect 28340 29892 28396 29894
rect 28420 29892 28476 29894
rect 28500 29892 28556 29894
rect 16180 21242 16236 21244
rect 16260 21242 16316 21244
rect 16340 21242 16396 21244
rect 16420 21242 16476 21244
rect 16500 21242 16556 21244
rect 16180 21190 16182 21242
rect 16182 21190 16234 21242
rect 16234 21190 16236 21242
rect 16260 21190 16298 21242
rect 16298 21190 16310 21242
rect 16310 21190 16316 21242
rect 16340 21190 16362 21242
rect 16362 21190 16374 21242
rect 16374 21190 16396 21242
rect 16420 21190 16426 21242
rect 16426 21190 16438 21242
rect 16438 21190 16476 21242
rect 16500 21190 16502 21242
rect 16502 21190 16554 21242
rect 16554 21190 16556 21242
rect 16180 21188 16236 21190
rect 16260 21188 16316 21190
rect 16340 21188 16396 21190
rect 16420 21188 16476 21190
rect 16500 21188 16556 21190
rect 16920 20698 16976 20700
rect 17000 20698 17056 20700
rect 17080 20698 17136 20700
rect 17160 20698 17216 20700
rect 17240 20698 17296 20700
rect 16920 20646 16922 20698
rect 16922 20646 16974 20698
rect 16974 20646 16976 20698
rect 17000 20646 17038 20698
rect 17038 20646 17050 20698
rect 17050 20646 17056 20698
rect 17080 20646 17102 20698
rect 17102 20646 17114 20698
rect 17114 20646 17136 20698
rect 17160 20646 17166 20698
rect 17166 20646 17178 20698
rect 17178 20646 17216 20698
rect 17240 20646 17242 20698
rect 17242 20646 17294 20698
rect 17294 20646 17296 20698
rect 16920 20644 16976 20646
rect 17000 20644 17056 20646
rect 17080 20644 17136 20646
rect 17160 20644 17216 20646
rect 17240 20644 17296 20646
rect 16180 20154 16236 20156
rect 16260 20154 16316 20156
rect 16340 20154 16396 20156
rect 16420 20154 16476 20156
rect 16500 20154 16556 20156
rect 16180 20102 16182 20154
rect 16182 20102 16234 20154
rect 16234 20102 16236 20154
rect 16260 20102 16298 20154
rect 16298 20102 16310 20154
rect 16310 20102 16316 20154
rect 16340 20102 16362 20154
rect 16362 20102 16374 20154
rect 16374 20102 16396 20154
rect 16420 20102 16426 20154
rect 16426 20102 16438 20154
rect 16438 20102 16476 20154
rect 16500 20102 16502 20154
rect 16502 20102 16554 20154
rect 16554 20102 16556 20154
rect 16180 20100 16236 20102
rect 16260 20100 16316 20102
rect 16340 20100 16396 20102
rect 16420 20100 16476 20102
rect 16500 20100 16556 20102
rect 16920 19610 16976 19612
rect 17000 19610 17056 19612
rect 17080 19610 17136 19612
rect 17160 19610 17216 19612
rect 17240 19610 17296 19612
rect 16920 19558 16922 19610
rect 16922 19558 16974 19610
rect 16974 19558 16976 19610
rect 17000 19558 17038 19610
rect 17038 19558 17050 19610
rect 17050 19558 17056 19610
rect 17080 19558 17102 19610
rect 17102 19558 17114 19610
rect 17114 19558 17136 19610
rect 17160 19558 17166 19610
rect 17166 19558 17178 19610
rect 17178 19558 17216 19610
rect 17240 19558 17242 19610
rect 17242 19558 17294 19610
rect 17294 19558 17296 19610
rect 16920 19556 16976 19558
rect 17000 19556 17056 19558
rect 17080 19556 17136 19558
rect 17160 19556 17216 19558
rect 17240 19556 17296 19558
rect 16180 19066 16236 19068
rect 16260 19066 16316 19068
rect 16340 19066 16396 19068
rect 16420 19066 16476 19068
rect 16500 19066 16556 19068
rect 16180 19014 16182 19066
rect 16182 19014 16234 19066
rect 16234 19014 16236 19066
rect 16260 19014 16298 19066
rect 16298 19014 16310 19066
rect 16310 19014 16316 19066
rect 16340 19014 16362 19066
rect 16362 19014 16374 19066
rect 16374 19014 16396 19066
rect 16420 19014 16426 19066
rect 16426 19014 16438 19066
rect 16438 19014 16476 19066
rect 16500 19014 16502 19066
rect 16502 19014 16554 19066
rect 16554 19014 16556 19066
rect 16180 19012 16236 19014
rect 16260 19012 16316 19014
rect 16340 19012 16396 19014
rect 16420 19012 16476 19014
rect 16500 19012 16556 19014
rect 16920 18522 16976 18524
rect 17000 18522 17056 18524
rect 17080 18522 17136 18524
rect 17160 18522 17216 18524
rect 17240 18522 17296 18524
rect 16920 18470 16922 18522
rect 16922 18470 16974 18522
rect 16974 18470 16976 18522
rect 17000 18470 17038 18522
rect 17038 18470 17050 18522
rect 17050 18470 17056 18522
rect 17080 18470 17102 18522
rect 17102 18470 17114 18522
rect 17114 18470 17136 18522
rect 17160 18470 17166 18522
rect 17166 18470 17178 18522
rect 17178 18470 17216 18522
rect 17240 18470 17242 18522
rect 17242 18470 17294 18522
rect 17294 18470 17296 18522
rect 16920 18468 16976 18470
rect 17000 18468 17056 18470
rect 17080 18468 17136 18470
rect 17160 18468 17216 18470
rect 17240 18468 17296 18470
rect 10920 5466 10976 5468
rect 11000 5466 11056 5468
rect 11080 5466 11136 5468
rect 11160 5466 11216 5468
rect 11240 5466 11296 5468
rect 10920 5414 10922 5466
rect 10922 5414 10974 5466
rect 10974 5414 10976 5466
rect 11000 5414 11038 5466
rect 11038 5414 11050 5466
rect 11050 5414 11056 5466
rect 11080 5414 11102 5466
rect 11102 5414 11114 5466
rect 11114 5414 11136 5466
rect 11160 5414 11166 5466
rect 11166 5414 11178 5466
rect 11178 5414 11216 5466
rect 11240 5414 11242 5466
rect 11242 5414 11294 5466
rect 11294 5414 11296 5466
rect 10920 5412 10976 5414
rect 11000 5412 11056 5414
rect 11080 5412 11136 5414
rect 11160 5412 11216 5414
rect 11240 5412 11296 5414
rect 10180 3834 10236 3836
rect 10260 3834 10316 3836
rect 10340 3834 10396 3836
rect 10420 3834 10476 3836
rect 10500 3834 10556 3836
rect 10180 3782 10182 3834
rect 10182 3782 10234 3834
rect 10234 3782 10236 3834
rect 10260 3782 10298 3834
rect 10298 3782 10310 3834
rect 10310 3782 10316 3834
rect 10340 3782 10362 3834
rect 10362 3782 10374 3834
rect 10374 3782 10396 3834
rect 10420 3782 10426 3834
rect 10426 3782 10438 3834
rect 10438 3782 10476 3834
rect 10500 3782 10502 3834
rect 10502 3782 10554 3834
rect 10554 3782 10556 3834
rect 10180 3780 10236 3782
rect 10260 3780 10316 3782
rect 10340 3780 10396 3782
rect 10420 3780 10476 3782
rect 10500 3780 10556 3782
rect 10920 4378 10976 4380
rect 11000 4378 11056 4380
rect 11080 4378 11136 4380
rect 11160 4378 11216 4380
rect 11240 4378 11296 4380
rect 10920 4326 10922 4378
rect 10922 4326 10974 4378
rect 10974 4326 10976 4378
rect 11000 4326 11038 4378
rect 11038 4326 11050 4378
rect 11050 4326 11056 4378
rect 11080 4326 11102 4378
rect 11102 4326 11114 4378
rect 11114 4326 11136 4378
rect 11160 4326 11166 4378
rect 11166 4326 11178 4378
rect 11178 4326 11216 4378
rect 11240 4326 11242 4378
rect 11242 4326 11294 4378
rect 11294 4326 11296 4378
rect 10920 4324 10976 4326
rect 11000 4324 11056 4326
rect 11080 4324 11136 4326
rect 11160 4324 11216 4326
rect 11240 4324 11296 4326
rect 10920 3290 10976 3292
rect 11000 3290 11056 3292
rect 11080 3290 11136 3292
rect 11160 3290 11216 3292
rect 11240 3290 11296 3292
rect 10920 3238 10922 3290
rect 10922 3238 10974 3290
rect 10974 3238 10976 3290
rect 11000 3238 11038 3290
rect 11038 3238 11050 3290
rect 11050 3238 11056 3290
rect 11080 3238 11102 3290
rect 11102 3238 11114 3290
rect 11114 3238 11136 3290
rect 11160 3238 11166 3290
rect 11166 3238 11178 3290
rect 11178 3238 11216 3290
rect 11240 3238 11242 3290
rect 11242 3238 11294 3290
rect 11294 3238 11296 3290
rect 10920 3236 10976 3238
rect 11000 3236 11056 3238
rect 11080 3236 11136 3238
rect 11160 3236 11216 3238
rect 11240 3236 11296 3238
rect 16180 17978 16236 17980
rect 16260 17978 16316 17980
rect 16340 17978 16396 17980
rect 16420 17978 16476 17980
rect 16500 17978 16556 17980
rect 16180 17926 16182 17978
rect 16182 17926 16234 17978
rect 16234 17926 16236 17978
rect 16260 17926 16298 17978
rect 16298 17926 16310 17978
rect 16310 17926 16316 17978
rect 16340 17926 16362 17978
rect 16362 17926 16374 17978
rect 16374 17926 16396 17978
rect 16420 17926 16426 17978
rect 16426 17926 16438 17978
rect 16438 17926 16476 17978
rect 16500 17926 16502 17978
rect 16502 17926 16554 17978
rect 16554 17926 16556 17978
rect 16180 17924 16236 17926
rect 16260 17924 16316 17926
rect 16340 17924 16396 17926
rect 16420 17924 16476 17926
rect 16500 17924 16556 17926
rect 16920 17434 16976 17436
rect 17000 17434 17056 17436
rect 17080 17434 17136 17436
rect 17160 17434 17216 17436
rect 17240 17434 17296 17436
rect 16920 17382 16922 17434
rect 16922 17382 16974 17434
rect 16974 17382 16976 17434
rect 17000 17382 17038 17434
rect 17038 17382 17050 17434
rect 17050 17382 17056 17434
rect 17080 17382 17102 17434
rect 17102 17382 17114 17434
rect 17114 17382 17136 17434
rect 17160 17382 17166 17434
rect 17166 17382 17178 17434
rect 17178 17382 17216 17434
rect 17240 17382 17242 17434
rect 17242 17382 17294 17434
rect 17294 17382 17296 17434
rect 16920 17380 16976 17382
rect 17000 17380 17056 17382
rect 17080 17380 17136 17382
rect 17160 17380 17216 17382
rect 17240 17380 17296 17382
rect 17866 17484 17868 17504
rect 17868 17484 17920 17504
rect 17920 17484 17922 17504
rect 17866 17448 17922 17484
rect 16180 16890 16236 16892
rect 16260 16890 16316 16892
rect 16340 16890 16396 16892
rect 16420 16890 16476 16892
rect 16500 16890 16556 16892
rect 16180 16838 16182 16890
rect 16182 16838 16234 16890
rect 16234 16838 16236 16890
rect 16260 16838 16298 16890
rect 16298 16838 16310 16890
rect 16310 16838 16316 16890
rect 16340 16838 16362 16890
rect 16362 16838 16374 16890
rect 16374 16838 16396 16890
rect 16420 16838 16426 16890
rect 16426 16838 16438 16890
rect 16438 16838 16476 16890
rect 16500 16838 16502 16890
rect 16502 16838 16554 16890
rect 16554 16838 16556 16890
rect 16180 16836 16236 16838
rect 16260 16836 16316 16838
rect 16340 16836 16396 16838
rect 16420 16836 16476 16838
rect 16500 16836 16556 16838
rect 16920 16346 16976 16348
rect 17000 16346 17056 16348
rect 17080 16346 17136 16348
rect 17160 16346 17216 16348
rect 17240 16346 17296 16348
rect 16920 16294 16922 16346
rect 16922 16294 16974 16346
rect 16974 16294 16976 16346
rect 17000 16294 17038 16346
rect 17038 16294 17050 16346
rect 17050 16294 17056 16346
rect 17080 16294 17102 16346
rect 17102 16294 17114 16346
rect 17114 16294 17136 16346
rect 17160 16294 17166 16346
rect 17166 16294 17178 16346
rect 17178 16294 17216 16346
rect 17240 16294 17242 16346
rect 17242 16294 17294 16346
rect 17294 16294 17296 16346
rect 16920 16292 16976 16294
rect 17000 16292 17056 16294
rect 17080 16292 17136 16294
rect 17160 16292 17216 16294
rect 17240 16292 17296 16294
rect 14830 8492 14886 8528
rect 18418 17604 18474 17640
rect 18418 17584 18420 17604
rect 18420 17584 18472 17604
rect 18472 17584 18474 17604
rect 16180 15802 16236 15804
rect 16260 15802 16316 15804
rect 16340 15802 16396 15804
rect 16420 15802 16476 15804
rect 16500 15802 16556 15804
rect 16180 15750 16182 15802
rect 16182 15750 16234 15802
rect 16234 15750 16236 15802
rect 16260 15750 16298 15802
rect 16298 15750 16310 15802
rect 16310 15750 16316 15802
rect 16340 15750 16362 15802
rect 16362 15750 16374 15802
rect 16374 15750 16396 15802
rect 16420 15750 16426 15802
rect 16426 15750 16438 15802
rect 16438 15750 16476 15802
rect 16500 15750 16502 15802
rect 16502 15750 16554 15802
rect 16554 15750 16556 15802
rect 16180 15748 16236 15750
rect 16260 15748 16316 15750
rect 16340 15748 16396 15750
rect 16420 15748 16476 15750
rect 16500 15748 16556 15750
rect 16920 15258 16976 15260
rect 17000 15258 17056 15260
rect 17080 15258 17136 15260
rect 17160 15258 17216 15260
rect 17240 15258 17296 15260
rect 16920 15206 16922 15258
rect 16922 15206 16974 15258
rect 16974 15206 16976 15258
rect 17000 15206 17038 15258
rect 17038 15206 17050 15258
rect 17050 15206 17056 15258
rect 17080 15206 17102 15258
rect 17102 15206 17114 15258
rect 17114 15206 17136 15258
rect 17160 15206 17166 15258
rect 17166 15206 17178 15258
rect 17178 15206 17216 15258
rect 17240 15206 17242 15258
rect 17242 15206 17294 15258
rect 17294 15206 17296 15258
rect 16920 15204 16976 15206
rect 17000 15204 17056 15206
rect 17080 15204 17136 15206
rect 17160 15204 17216 15206
rect 17240 15204 17296 15206
rect 16180 14714 16236 14716
rect 16260 14714 16316 14716
rect 16340 14714 16396 14716
rect 16420 14714 16476 14716
rect 16500 14714 16556 14716
rect 16180 14662 16182 14714
rect 16182 14662 16234 14714
rect 16234 14662 16236 14714
rect 16260 14662 16298 14714
rect 16298 14662 16310 14714
rect 16310 14662 16316 14714
rect 16340 14662 16362 14714
rect 16362 14662 16374 14714
rect 16374 14662 16396 14714
rect 16420 14662 16426 14714
rect 16426 14662 16438 14714
rect 16438 14662 16476 14714
rect 16500 14662 16502 14714
rect 16502 14662 16554 14714
rect 16554 14662 16556 14714
rect 16180 14660 16236 14662
rect 16260 14660 16316 14662
rect 16340 14660 16396 14662
rect 16420 14660 16476 14662
rect 16500 14660 16556 14662
rect 16920 14170 16976 14172
rect 17000 14170 17056 14172
rect 17080 14170 17136 14172
rect 17160 14170 17216 14172
rect 17240 14170 17296 14172
rect 16920 14118 16922 14170
rect 16922 14118 16974 14170
rect 16974 14118 16976 14170
rect 17000 14118 17038 14170
rect 17038 14118 17050 14170
rect 17050 14118 17056 14170
rect 17080 14118 17102 14170
rect 17102 14118 17114 14170
rect 17114 14118 17136 14170
rect 17160 14118 17166 14170
rect 17166 14118 17178 14170
rect 17178 14118 17216 14170
rect 17240 14118 17242 14170
rect 17242 14118 17294 14170
rect 17294 14118 17296 14170
rect 16920 14116 16976 14118
rect 17000 14116 17056 14118
rect 17080 14116 17136 14118
rect 17160 14116 17216 14118
rect 17240 14116 17296 14118
rect 14830 8472 14832 8492
rect 14832 8472 14884 8492
rect 14884 8472 14886 8492
rect 15382 7248 15438 7304
rect 16180 13626 16236 13628
rect 16260 13626 16316 13628
rect 16340 13626 16396 13628
rect 16420 13626 16476 13628
rect 16500 13626 16556 13628
rect 16180 13574 16182 13626
rect 16182 13574 16234 13626
rect 16234 13574 16236 13626
rect 16260 13574 16298 13626
rect 16298 13574 16310 13626
rect 16310 13574 16316 13626
rect 16340 13574 16362 13626
rect 16362 13574 16374 13626
rect 16374 13574 16396 13626
rect 16420 13574 16426 13626
rect 16426 13574 16438 13626
rect 16438 13574 16476 13626
rect 16500 13574 16502 13626
rect 16502 13574 16554 13626
rect 16554 13574 16556 13626
rect 16180 13572 16236 13574
rect 16260 13572 16316 13574
rect 16340 13572 16396 13574
rect 16420 13572 16476 13574
rect 16500 13572 16556 13574
rect 16920 13082 16976 13084
rect 17000 13082 17056 13084
rect 17080 13082 17136 13084
rect 17160 13082 17216 13084
rect 17240 13082 17296 13084
rect 16920 13030 16922 13082
rect 16922 13030 16974 13082
rect 16974 13030 16976 13082
rect 17000 13030 17038 13082
rect 17038 13030 17050 13082
rect 17050 13030 17056 13082
rect 17080 13030 17102 13082
rect 17102 13030 17114 13082
rect 17114 13030 17136 13082
rect 17160 13030 17166 13082
rect 17166 13030 17178 13082
rect 17178 13030 17216 13082
rect 17240 13030 17242 13082
rect 17242 13030 17294 13082
rect 17294 13030 17296 13082
rect 16920 13028 16976 13030
rect 17000 13028 17056 13030
rect 17080 13028 17136 13030
rect 17160 13028 17216 13030
rect 17240 13028 17296 13030
rect 16180 12538 16236 12540
rect 16260 12538 16316 12540
rect 16340 12538 16396 12540
rect 16420 12538 16476 12540
rect 16500 12538 16556 12540
rect 16180 12486 16182 12538
rect 16182 12486 16234 12538
rect 16234 12486 16236 12538
rect 16260 12486 16298 12538
rect 16298 12486 16310 12538
rect 16310 12486 16316 12538
rect 16340 12486 16362 12538
rect 16362 12486 16374 12538
rect 16374 12486 16396 12538
rect 16420 12486 16426 12538
rect 16426 12486 16438 12538
rect 16438 12486 16476 12538
rect 16500 12486 16502 12538
rect 16502 12486 16554 12538
rect 16554 12486 16556 12538
rect 16180 12484 16236 12486
rect 16260 12484 16316 12486
rect 16340 12484 16396 12486
rect 16420 12484 16476 12486
rect 16500 12484 16556 12486
rect 16920 11994 16976 11996
rect 17000 11994 17056 11996
rect 17080 11994 17136 11996
rect 17160 11994 17216 11996
rect 17240 11994 17296 11996
rect 16920 11942 16922 11994
rect 16922 11942 16974 11994
rect 16974 11942 16976 11994
rect 17000 11942 17038 11994
rect 17038 11942 17050 11994
rect 17050 11942 17056 11994
rect 17080 11942 17102 11994
rect 17102 11942 17114 11994
rect 17114 11942 17136 11994
rect 17160 11942 17166 11994
rect 17166 11942 17178 11994
rect 17178 11942 17216 11994
rect 17240 11942 17242 11994
rect 17242 11942 17294 11994
rect 17294 11942 17296 11994
rect 16920 11940 16976 11942
rect 17000 11940 17056 11942
rect 17080 11940 17136 11942
rect 17160 11940 17216 11942
rect 17240 11940 17296 11942
rect 16180 11450 16236 11452
rect 16260 11450 16316 11452
rect 16340 11450 16396 11452
rect 16420 11450 16476 11452
rect 16500 11450 16556 11452
rect 16180 11398 16182 11450
rect 16182 11398 16234 11450
rect 16234 11398 16236 11450
rect 16260 11398 16298 11450
rect 16298 11398 16310 11450
rect 16310 11398 16316 11450
rect 16340 11398 16362 11450
rect 16362 11398 16374 11450
rect 16374 11398 16396 11450
rect 16420 11398 16426 11450
rect 16426 11398 16438 11450
rect 16438 11398 16476 11450
rect 16500 11398 16502 11450
rect 16502 11398 16554 11450
rect 16554 11398 16556 11450
rect 16180 11396 16236 11398
rect 16260 11396 16316 11398
rect 16340 11396 16396 11398
rect 16420 11396 16476 11398
rect 16500 11396 16556 11398
rect 16920 10906 16976 10908
rect 17000 10906 17056 10908
rect 17080 10906 17136 10908
rect 17160 10906 17216 10908
rect 17240 10906 17296 10908
rect 16920 10854 16922 10906
rect 16922 10854 16974 10906
rect 16974 10854 16976 10906
rect 17000 10854 17038 10906
rect 17038 10854 17050 10906
rect 17050 10854 17056 10906
rect 17080 10854 17102 10906
rect 17102 10854 17114 10906
rect 17114 10854 17136 10906
rect 17160 10854 17166 10906
rect 17166 10854 17178 10906
rect 17178 10854 17216 10906
rect 17240 10854 17242 10906
rect 17242 10854 17294 10906
rect 17294 10854 17296 10906
rect 16920 10852 16976 10854
rect 17000 10852 17056 10854
rect 17080 10852 17136 10854
rect 17160 10852 17216 10854
rect 17240 10852 17296 10854
rect 16180 10362 16236 10364
rect 16260 10362 16316 10364
rect 16340 10362 16396 10364
rect 16420 10362 16476 10364
rect 16500 10362 16556 10364
rect 16180 10310 16182 10362
rect 16182 10310 16234 10362
rect 16234 10310 16236 10362
rect 16260 10310 16298 10362
rect 16298 10310 16310 10362
rect 16310 10310 16316 10362
rect 16340 10310 16362 10362
rect 16362 10310 16374 10362
rect 16374 10310 16396 10362
rect 16420 10310 16426 10362
rect 16426 10310 16438 10362
rect 16438 10310 16476 10362
rect 16500 10310 16502 10362
rect 16502 10310 16554 10362
rect 16554 10310 16556 10362
rect 16180 10308 16236 10310
rect 16260 10308 16316 10310
rect 16340 10308 16396 10310
rect 16420 10308 16476 10310
rect 16500 10308 16556 10310
rect 16920 9818 16976 9820
rect 17000 9818 17056 9820
rect 17080 9818 17136 9820
rect 17160 9818 17216 9820
rect 17240 9818 17296 9820
rect 16920 9766 16922 9818
rect 16922 9766 16974 9818
rect 16974 9766 16976 9818
rect 17000 9766 17038 9818
rect 17038 9766 17050 9818
rect 17050 9766 17056 9818
rect 17080 9766 17102 9818
rect 17102 9766 17114 9818
rect 17114 9766 17136 9818
rect 17160 9766 17166 9818
rect 17166 9766 17178 9818
rect 17178 9766 17216 9818
rect 17240 9766 17242 9818
rect 17242 9766 17294 9818
rect 17294 9766 17296 9818
rect 16920 9764 16976 9766
rect 17000 9764 17056 9766
rect 17080 9764 17136 9766
rect 17160 9764 17216 9766
rect 17240 9764 17296 9766
rect 16180 9274 16236 9276
rect 16260 9274 16316 9276
rect 16340 9274 16396 9276
rect 16420 9274 16476 9276
rect 16500 9274 16556 9276
rect 16180 9222 16182 9274
rect 16182 9222 16234 9274
rect 16234 9222 16236 9274
rect 16260 9222 16298 9274
rect 16298 9222 16310 9274
rect 16310 9222 16316 9274
rect 16340 9222 16362 9274
rect 16362 9222 16374 9274
rect 16374 9222 16396 9274
rect 16420 9222 16426 9274
rect 16426 9222 16438 9274
rect 16438 9222 16476 9274
rect 16500 9222 16502 9274
rect 16502 9222 16554 9274
rect 16554 9222 16556 9274
rect 16180 9220 16236 9222
rect 16260 9220 16316 9222
rect 16340 9220 16396 9222
rect 16420 9220 16476 9222
rect 16500 9220 16556 9222
rect 16920 8730 16976 8732
rect 17000 8730 17056 8732
rect 17080 8730 17136 8732
rect 17160 8730 17216 8732
rect 17240 8730 17296 8732
rect 16920 8678 16922 8730
rect 16922 8678 16974 8730
rect 16974 8678 16976 8730
rect 17000 8678 17038 8730
rect 17038 8678 17050 8730
rect 17050 8678 17056 8730
rect 17080 8678 17102 8730
rect 17102 8678 17114 8730
rect 17114 8678 17136 8730
rect 17160 8678 17166 8730
rect 17166 8678 17178 8730
rect 17178 8678 17216 8730
rect 17240 8678 17242 8730
rect 17242 8678 17294 8730
rect 17294 8678 17296 8730
rect 16920 8676 16976 8678
rect 17000 8676 17056 8678
rect 17080 8676 17136 8678
rect 17160 8676 17216 8678
rect 17240 8676 17296 8678
rect 16180 8186 16236 8188
rect 16260 8186 16316 8188
rect 16340 8186 16396 8188
rect 16420 8186 16476 8188
rect 16500 8186 16556 8188
rect 16180 8134 16182 8186
rect 16182 8134 16234 8186
rect 16234 8134 16236 8186
rect 16260 8134 16298 8186
rect 16298 8134 16310 8186
rect 16310 8134 16316 8186
rect 16340 8134 16362 8186
rect 16362 8134 16374 8186
rect 16374 8134 16396 8186
rect 16420 8134 16426 8186
rect 16426 8134 16438 8186
rect 16438 8134 16476 8186
rect 16500 8134 16502 8186
rect 16502 8134 16554 8186
rect 16554 8134 16556 8186
rect 16180 8132 16236 8134
rect 16260 8132 16316 8134
rect 16340 8132 16396 8134
rect 16420 8132 16476 8134
rect 16500 8132 16556 8134
rect 16180 7098 16236 7100
rect 16260 7098 16316 7100
rect 16340 7098 16396 7100
rect 16420 7098 16476 7100
rect 16500 7098 16556 7100
rect 16180 7046 16182 7098
rect 16182 7046 16234 7098
rect 16234 7046 16236 7098
rect 16260 7046 16298 7098
rect 16298 7046 16310 7098
rect 16310 7046 16316 7098
rect 16340 7046 16362 7098
rect 16362 7046 16374 7098
rect 16374 7046 16396 7098
rect 16420 7046 16426 7098
rect 16426 7046 16438 7098
rect 16438 7046 16476 7098
rect 16500 7046 16502 7098
rect 16502 7046 16554 7098
rect 16554 7046 16556 7098
rect 16180 7044 16236 7046
rect 16260 7044 16316 7046
rect 16340 7044 16396 7046
rect 16420 7044 16476 7046
rect 16500 7044 16556 7046
rect 16920 7642 16976 7644
rect 17000 7642 17056 7644
rect 17080 7642 17136 7644
rect 17160 7642 17216 7644
rect 17240 7642 17296 7644
rect 16920 7590 16922 7642
rect 16922 7590 16974 7642
rect 16974 7590 16976 7642
rect 17000 7590 17038 7642
rect 17038 7590 17050 7642
rect 17050 7590 17056 7642
rect 17080 7590 17102 7642
rect 17102 7590 17114 7642
rect 17114 7590 17136 7642
rect 17160 7590 17166 7642
rect 17166 7590 17178 7642
rect 17178 7590 17216 7642
rect 17240 7590 17242 7642
rect 17242 7590 17294 7642
rect 17294 7590 17296 7642
rect 16920 7588 16976 7590
rect 17000 7588 17056 7590
rect 17080 7588 17136 7590
rect 17160 7588 17216 7590
rect 17240 7588 17296 7590
rect 16180 6010 16236 6012
rect 16260 6010 16316 6012
rect 16340 6010 16396 6012
rect 16420 6010 16476 6012
rect 16500 6010 16556 6012
rect 16180 5958 16182 6010
rect 16182 5958 16234 6010
rect 16234 5958 16236 6010
rect 16260 5958 16298 6010
rect 16298 5958 16310 6010
rect 16310 5958 16316 6010
rect 16340 5958 16362 6010
rect 16362 5958 16374 6010
rect 16374 5958 16396 6010
rect 16420 5958 16426 6010
rect 16426 5958 16438 6010
rect 16438 5958 16476 6010
rect 16500 5958 16502 6010
rect 16502 5958 16554 6010
rect 16554 5958 16556 6010
rect 16180 5956 16236 5958
rect 16260 5956 16316 5958
rect 16340 5956 16396 5958
rect 16420 5956 16476 5958
rect 16500 5956 16556 5958
rect 17314 6704 17370 6760
rect 16920 6554 16976 6556
rect 17000 6554 17056 6556
rect 17080 6554 17136 6556
rect 17160 6554 17216 6556
rect 17240 6554 17296 6556
rect 16920 6502 16922 6554
rect 16922 6502 16974 6554
rect 16974 6502 16976 6554
rect 17000 6502 17038 6554
rect 17038 6502 17050 6554
rect 17050 6502 17056 6554
rect 17080 6502 17102 6554
rect 17102 6502 17114 6554
rect 17114 6502 17136 6554
rect 17160 6502 17166 6554
rect 17166 6502 17178 6554
rect 17178 6502 17216 6554
rect 17240 6502 17242 6554
rect 17242 6502 17294 6554
rect 17294 6502 17296 6554
rect 16920 6500 16976 6502
rect 17000 6500 17056 6502
rect 17080 6500 17136 6502
rect 17160 6500 17216 6502
rect 17240 6500 17296 6502
rect 22920 29402 22976 29404
rect 23000 29402 23056 29404
rect 23080 29402 23136 29404
rect 23160 29402 23216 29404
rect 23240 29402 23296 29404
rect 22920 29350 22922 29402
rect 22922 29350 22974 29402
rect 22974 29350 22976 29402
rect 23000 29350 23038 29402
rect 23038 29350 23050 29402
rect 23050 29350 23056 29402
rect 23080 29350 23102 29402
rect 23102 29350 23114 29402
rect 23114 29350 23136 29402
rect 23160 29350 23166 29402
rect 23166 29350 23178 29402
rect 23178 29350 23216 29402
rect 23240 29350 23242 29402
rect 23242 29350 23294 29402
rect 23294 29350 23296 29402
rect 22920 29348 22976 29350
rect 23000 29348 23056 29350
rect 23080 29348 23136 29350
rect 23160 29348 23216 29350
rect 23240 29348 23296 29350
rect 28920 29402 28976 29404
rect 29000 29402 29056 29404
rect 29080 29402 29136 29404
rect 29160 29402 29216 29404
rect 29240 29402 29296 29404
rect 28920 29350 28922 29402
rect 28922 29350 28974 29402
rect 28974 29350 28976 29402
rect 29000 29350 29038 29402
rect 29038 29350 29050 29402
rect 29050 29350 29056 29402
rect 29080 29350 29102 29402
rect 29102 29350 29114 29402
rect 29114 29350 29136 29402
rect 29160 29350 29166 29402
rect 29166 29350 29178 29402
rect 29178 29350 29216 29402
rect 29240 29350 29242 29402
rect 29242 29350 29294 29402
rect 29294 29350 29296 29402
rect 28920 29348 28976 29350
rect 29000 29348 29056 29350
rect 29080 29348 29136 29350
rect 29160 29348 29216 29350
rect 29240 29348 29296 29350
rect 22180 28858 22236 28860
rect 22260 28858 22316 28860
rect 22340 28858 22396 28860
rect 22420 28858 22476 28860
rect 22500 28858 22556 28860
rect 22180 28806 22182 28858
rect 22182 28806 22234 28858
rect 22234 28806 22236 28858
rect 22260 28806 22298 28858
rect 22298 28806 22310 28858
rect 22310 28806 22316 28858
rect 22340 28806 22362 28858
rect 22362 28806 22374 28858
rect 22374 28806 22396 28858
rect 22420 28806 22426 28858
rect 22426 28806 22438 28858
rect 22438 28806 22476 28858
rect 22500 28806 22502 28858
rect 22502 28806 22554 28858
rect 22554 28806 22556 28858
rect 22180 28804 22236 28806
rect 22260 28804 22316 28806
rect 22340 28804 22396 28806
rect 22420 28804 22476 28806
rect 22500 28804 22556 28806
rect 28180 28858 28236 28860
rect 28260 28858 28316 28860
rect 28340 28858 28396 28860
rect 28420 28858 28476 28860
rect 28500 28858 28556 28860
rect 28180 28806 28182 28858
rect 28182 28806 28234 28858
rect 28234 28806 28236 28858
rect 28260 28806 28298 28858
rect 28298 28806 28310 28858
rect 28310 28806 28316 28858
rect 28340 28806 28362 28858
rect 28362 28806 28374 28858
rect 28374 28806 28396 28858
rect 28420 28806 28426 28858
rect 28426 28806 28438 28858
rect 28438 28806 28476 28858
rect 28500 28806 28502 28858
rect 28502 28806 28554 28858
rect 28554 28806 28556 28858
rect 28180 28804 28236 28806
rect 28260 28804 28316 28806
rect 28340 28804 28396 28806
rect 28420 28804 28476 28806
rect 28500 28804 28556 28806
rect 22920 28314 22976 28316
rect 23000 28314 23056 28316
rect 23080 28314 23136 28316
rect 23160 28314 23216 28316
rect 23240 28314 23296 28316
rect 22920 28262 22922 28314
rect 22922 28262 22974 28314
rect 22974 28262 22976 28314
rect 23000 28262 23038 28314
rect 23038 28262 23050 28314
rect 23050 28262 23056 28314
rect 23080 28262 23102 28314
rect 23102 28262 23114 28314
rect 23114 28262 23136 28314
rect 23160 28262 23166 28314
rect 23166 28262 23178 28314
rect 23178 28262 23216 28314
rect 23240 28262 23242 28314
rect 23242 28262 23294 28314
rect 23294 28262 23296 28314
rect 22920 28260 22976 28262
rect 23000 28260 23056 28262
rect 23080 28260 23136 28262
rect 23160 28260 23216 28262
rect 23240 28260 23296 28262
rect 28920 28314 28976 28316
rect 29000 28314 29056 28316
rect 29080 28314 29136 28316
rect 29160 28314 29216 28316
rect 29240 28314 29296 28316
rect 28920 28262 28922 28314
rect 28922 28262 28974 28314
rect 28974 28262 28976 28314
rect 29000 28262 29038 28314
rect 29038 28262 29050 28314
rect 29050 28262 29056 28314
rect 29080 28262 29102 28314
rect 29102 28262 29114 28314
rect 29114 28262 29136 28314
rect 29160 28262 29166 28314
rect 29166 28262 29178 28314
rect 29178 28262 29216 28314
rect 29240 28262 29242 28314
rect 29242 28262 29294 28314
rect 29294 28262 29296 28314
rect 28920 28260 28976 28262
rect 29000 28260 29056 28262
rect 29080 28260 29136 28262
rect 29160 28260 29216 28262
rect 29240 28260 29296 28262
rect 22180 27770 22236 27772
rect 22260 27770 22316 27772
rect 22340 27770 22396 27772
rect 22420 27770 22476 27772
rect 22500 27770 22556 27772
rect 22180 27718 22182 27770
rect 22182 27718 22234 27770
rect 22234 27718 22236 27770
rect 22260 27718 22298 27770
rect 22298 27718 22310 27770
rect 22310 27718 22316 27770
rect 22340 27718 22362 27770
rect 22362 27718 22374 27770
rect 22374 27718 22396 27770
rect 22420 27718 22426 27770
rect 22426 27718 22438 27770
rect 22438 27718 22476 27770
rect 22500 27718 22502 27770
rect 22502 27718 22554 27770
rect 22554 27718 22556 27770
rect 22180 27716 22236 27718
rect 22260 27716 22316 27718
rect 22340 27716 22396 27718
rect 22420 27716 22476 27718
rect 22500 27716 22556 27718
rect 22180 26682 22236 26684
rect 22260 26682 22316 26684
rect 22340 26682 22396 26684
rect 22420 26682 22476 26684
rect 22500 26682 22556 26684
rect 22180 26630 22182 26682
rect 22182 26630 22234 26682
rect 22234 26630 22236 26682
rect 22260 26630 22298 26682
rect 22298 26630 22310 26682
rect 22310 26630 22316 26682
rect 22340 26630 22362 26682
rect 22362 26630 22374 26682
rect 22374 26630 22396 26682
rect 22420 26630 22426 26682
rect 22426 26630 22438 26682
rect 22438 26630 22476 26682
rect 22500 26630 22502 26682
rect 22502 26630 22554 26682
rect 22554 26630 22556 26682
rect 22180 26628 22236 26630
rect 22260 26628 22316 26630
rect 22340 26628 22396 26630
rect 22420 26628 22476 26630
rect 22500 26628 22556 26630
rect 20718 21528 20774 21584
rect 20718 20712 20774 20768
rect 22920 27226 22976 27228
rect 23000 27226 23056 27228
rect 23080 27226 23136 27228
rect 23160 27226 23216 27228
rect 23240 27226 23296 27228
rect 22920 27174 22922 27226
rect 22922 27174 22974 27226
rect 22974 27174 22976 27226
rect 23000 27174 23038 27226
rect 23038 27174 23050 27226
rect 23050 27174 23056 27226
rect 23080 27174 23102 27226
rect 23102 27174 23114 27226
rect 23114 27174 23136 27226
rect 23160 27174 23166 27226
rect 23166 27174 23178 27226
rect 23178 27174 23216 27226
rect 23240 27174 23242 27226
rect 23242 27174 23294 27226
rect 23294 27174 23296 27226
rect 22920 27172 22976 27174
rect 23000 27172 23056 27174
rect 23080 27172 23136 27174
rect 23160 27172 23216 27174
rect 23240 27172 23296 27174
rect 23754 26988 23810 27024
rect 23754 26968 23756 26988
rect 23756 26968 23808 26988
rect 23808 26968 23810 26988
rect 22920 26138 22976 26140
rect 23000 26138 23056 26140
rect 23080 26138 23136 26140
rect 23160 26138 23216 26140
rect 23240 26138 23296 26140
rect 22920 26086 22922 26138
rect 22922 26086 22974 26138
rect 22974 26086 22976 26138
rect 23000 26086 23038 26138
rect 23038 26086 23050 26138
rect 23050 26086 23056 26138
rect 23080 26086 23102 26138
rect 23102 26086 23114 26138
rect 23114 26086 23136 26138
rect 23160 26086 23166 26138
rect 23166 26086 23178 26138
rect 23178 26086 23216 26138
rect 23240 26086 23242 26138
rect 23242 26086 23294 26138
rect 23294 26086 23296 26138
rect 22920 26084 22976 26086
rect 23000 26084 23056 26086
rect 23080 26084 23136 26086
rect 23160 26084 23216 26086
rect 23240 26084 23296 26086
rect 22180 25594 22236 25596
rect 22260 25594 22316 25596
rect 22340 25594 22396 25596
rect 22420 25594 22476 25596
rect 22500 25594 22556 25596
rect 22180 25542 22182 25594
rect 22182 25542 22234 25594
rect 22234 25542 22236 25594
rect 22260 25542 22298 25594
rect 22298 25542 22310 25594
rect 22310 25542 22316 25594
rect 22340 25542 22362 25594
rect 22362 25542 22374 25594
rect 22374 25542 22396 25594
rect 22420 25542 22426 25594
rect 22426 25542 22438 25594
rect 22438 25542 22476 25594
rect 22500 25542 22502 25594
rect 22502 25542 22554 25594
rect 22554 25542 22556 25594
rect 22180 25540 22236 25542
rect 22260 25540 22316 25542
rect 22340 25540 22396 25542
rect 22420 25540 22476 25542
rect 22500 25540 22556 25542
rect 22920 25050 22976 25052
rect 23000 25050 23056 25052
rect 23080 25050 23136 25052
rect 23160 25050 23216 25052
rect 23240 25050 23296 25052
rect 22920 24998 22922 25050
rect 22922 24998 22974 25050
rect 22974 24998 22976 25050
rect 23000 24998 23038 25050
rect 23038 24998 23050 25050
rect 23050 24998 23056 25050
rect 23080 24998 23102 25050
rect 23102 24998 23114 25050
rect 23114 24998 23136 25050
rect 23160 24998 23166 25050
rect 23166 24998 23178 25050
rect 23178 24998 23216 25050
rect 23240 24998 23242 25050
rect 23242 24998 23294 25050
rect 23294 24998 23296 25050
rect 22920 24996 22976 24998
rect 23000 24996 23056 24998
rect 23080 24996 23136 24998
rect 23160 24996 23216 24998
rect 23240 24996 23296 24998
rect 22180 24506 22236 24508
rect 22260 24506 22316 24508
rect 22340 24506 22396 24508
rect 22420 24506 22476 24508
rect 22500 24506 22556 24508
rect 22180 24454 22182 24506
rect 22182 24454 22234 24506
rect 22234 24454 22236 24506
rect 22260 24454 22298 24506
rect 22298 24454 22310 24506
rect 22310 24454 22316 24506
rect 22340 24454 22362 24506
rect 22362 24454 22374 24506
rect 22374 24454 22396 24506
rect 22420 24454 22426 24506
rect 22426 24454 22438 24506
rect 22438 24454 22476 24506
rect 22500 24454 22502 24506
rect 22502 24454 22554 24506
rect 22554 24454 22556 24506
rect 22180 24452 22236 24454
rect 22260 24452 22316 24454
rect 22340 24452 22396 24454
rect 22420 24452 22476 24454
rect 22500 24452 22556 24454
rect 22920 23962 22976 23964
rect 23000 23962 23056 23964
rect 23080 23962 23136 23964
rect 23160 23962 23216 23964
rect 23240 23962 23296 23964
rect 22920 23910 22922 23962
rect 22922 23910 22974 23962
rect 22974 23910 22976 23962
rect 23000 23910 23038 23962
rect 23038 23910 23050 23962
rect 23050 23910 23056 23962
rect 23080 23910 23102 23962
rect 23102 23910 23114 23962
rect 23114 23910 23136 23962
rect 23160 23910 23166 23962
rect 23166 23910 23178 23962
rect 23178 23910 23216 23962
rect 23240 23910 23242 23962
rect 23242 23910 23294 23962
rect 23294 23910 23296 23962
rect 22920 23908 22976 23910
rect 23000 23908 23056 23910
rect 23080 23908 23136 23910
rect 23160 23908 23216 23910
rect 23240 23908 23296 23910
rect 22180 23418 22236 23420
rect 22260 23418 22316 23420
rect 22340 23418 22396 23420
rect 22420 23418 22476 23420
rect 22500 23418 22556 23420
rect 22180 23366 22182 23418
rect 22182 23366 22234 23418
rect 22234 23366 22236 23418
rect 22260 23366 22298 23418
rect 22298 23366 22310 23418
rect 22310 23366 22316 23418
rect 22340 23366 22362 23418
rect 22362 23366 22374 23418
rect 22374 23366 22396 23418
rect 22420 23366 22426 23418
rect 22426 23366 22438 23418
rect 22438 23366 22476 23418
rect 22500 23366 22502 23418
rect 22502 23366 22554 23418
rect 22554 23366 22556 23418
rect 22180 23364 22236 23366
rect 22260 23364 22316 23366
rect 22340 23364 22396 23366
rect 22420 23364 22476 23366
rect 22500 23364 22556 23366
rect 22180 22330 22236 22332
rect 22260 22330 22316 22332
rect 22340 22330 22396 22332
rect 22420 22330 22476 22332
rect 22500 22330 22556 22332
rect 22180 22278 22182 22330
rect 22182 22278 22234 22330
rect 22234 22278 22236 22330
rect 22260 22278 22298 22330
rect 22298 22278 22310 22330
rect 22310 22278 22316 22330
rect 22340 22278 22362 22330
rect 22362 22278 22374 22330
rect 22374 22278 22396 22330
rect 22420 22278 22426 22330
rect 22426 22278 22438 22330
rect 22438 22278 22476 22330
rect 22500 22278 22502 22330
rect 22502 22278 22554 22330
rect 22554 22278 22556 22330
rect 22180 22276 22236 22278
rect 22260 22276 22316 22278
rect 22340 22276 22396 22278
rect 22420 22276 22476 22278
rect 22500 22276 22556 22278
rect 22180 21242 22236 21244
rect 22260 21242 22316 21244
rect 22340 21242 22396 21244
rect 22420 21242 22476 21244
rect 22500 21242 22556 21244
rect 22180 21190 22182 21242
rect 22182 21190 22234 21242
rect 22234 21190 22236 21242
rect 22260 21190 22298 21242
rect 22298 21190 22310 21242
rect 22310 21190 22316 21242
rect 22340 21190 22362 21242
rect 22362 21190 22374 21242
rect 22374 21190 22396 21242
rect 22420 21190 22426 21242
rect 22426 21190 22438 21242
rect 22438 21190 22476 21242
rect 22500 21190 22502 21242
rect 22502 21190 22554 21242
rect 22554 21190 22556 21242
rect 22180 21188 22236 21190
rect 22260 21188 22316 21190
rect 22340 21188 22396 21190
rect 22420 21188 22476 21190
rect 22500 21188 22556 21190
rect 22180 20154 22236 20156
rect 22260 20154 22316 20156
rect 22340 20154 22396 20156
rect 22420 20154 22476 20156
rect 22500 20154 22556 20156
rect 22180 20102 22182 20154
rect 22182 20102 22234 20154
rect 22234 20102 22236 20154
rect 22260 20102 22298 20154
rect 22298 20102 22310 20154
rect 22310 20102 22316 20154
rect 22340 20102 22362 20154
rect 22362 20102 22374 20154
rect 22374 20102 22396 20154
rect 22420 20102 22426 20154
rect 22426 20102 22438 20154
rect 22438 20102 22476 20154
rect 22500 20102 22502 20154
rect 22502 20102 22554 20154
rect 22554 20102 22556 20154
rect 22180 20100 22236 20102
rect 22260 20100 22316 20102
rect 22340 20100 22396 20102
rect 22420 20100 22476 20102
rect 22500 20100 22556 20102
rect 22920 22874 22976 22876
rect 23000 22874 23056 22876
rect 23080 22874 23136 22876
rect 23160 22874 23216 22876
rect 23240 22874 23296 22876
rect 22920 22822 22922 22874
rect 22922 22822 22974 22874
rect 22974 22822 22976 22874
rect 23000 22822 23038 22874
rect 23038 22822 23050 22874
rect 23050 22822 23056 22874
rect 23080 22822 23102 22874
rect 23102 22822 23114 22874
rect 23114 22822 23136 22874
rect 23160 22822 23166 22874
rect 23166 22822 23178 22874
rect 23178 22822 23216 22874
rect 23240 22822 23242 22874
rect 23242 22822 23294 22874
rect 23294 22822 23296 22874
rect 22920 22820 22976 22822
rect 23000 22820 23056 22822
rect 23080 22820 23136 22822
rect 23160 22820 23216 22822
rect 23240 22820 23296 22822
rect 22920 21786 22976 21788
rect 23000 21786 23056 21788
rect 23080 21786 23136 21788
rect 23160 21786 23216 21788
rect 23240 21786 23296 21788
rect 22920 21734 22922 21786
rect 22922 21734 22974 21786
rect 22974 21734 22976 21786
rect 23000 21734 23038 21786
rect 23038 21734 23050 21786
rect 23050 21734 23056 21786
rect 23080 21734 23102 21786
rect 23102 21734 23114 21786
rect 23114 21734 23136 21786
rect 23160 21734 23166 21786
rect 23166 21734 23178 21786
rect 23178 21734 23216 21786
rect 23240 21734 23242 21786
rect 23242 21734 23294 21786
rect 23294 21734 23296 21786
rect 22920 21732 22976 21734
rect 23000 21732 23056 21734
rect 23080 21732 23136 21734
rect 23160 21732 23216 21734
rect 23240 21732 23296 21734
rect 22920 20698 22976 20700
rect 23000 20698 23056 20700
rect 23080 20698 23136 20700
rect 23160 20698 23216 20700
rect 23240 20698 23296 20700
rect 22920 20646 22922 20698
rect 22922 20646 22974 20698
rect 22974 20646 22976 20698
rect 23000 20646 23038 20698
rect 23038 20646 23050 20698
rect 23050 20646 23056 20698
rect 23080 20646 23102 20698
rect 23102 20646 23114 20698
rect 23114 20646 23136 20698
rect 23160 20646 23166 20698
rect 23166 20646 23178 20698
rect 23178 20646 23216 20698
rect 23240 20646 23242 20698
rect 23242 20646 23294 20698
rect 23294 20646 23296 20698
rect 22920 20644 22976 20646
rect 23000 20644 23056 20646
rect 23080 20644 23136 20646
rect 23160 20644 23216 20646
rect 23240 20644 23296 20646
rect 22180 19066 22236 19068
rect 22260 19066 22316 19068
rect 22340 19066 22396 19068
rect 22420 19066 22476 19068
rect 22500 19066 22556 19068
rect 22180 19014 22182 19066
rect 22182 19014 22234 19066
rect 22234 19014 22236 19066
rect 22260 19014 22298 19066
rect 22298 19014 22310 19066
rect 22310 19014 22316 19066
rect 22340 19014 22362 19066
rect 22362 19014 22374 19066
rect 22374 19014 22396 19066
rect 22420 19014 22426 19066
rect 22426 19014 22438 19066
rect 22438 19014 22476 19066
rect 22500 19014 22502 19066
rect 22502 19014 22554 19066
rect 22554 19014 22556 19066
rect 22180 19012 22236 19014
rect 22260 19012 22316 19014
rect 22340 19012 22396 19014
rect 22420 19012 22476 19014
rect 22500 19012 22556 19014
rect 22920 19610 22976 19612
rect 23000 19610 23056 19612
rect 23080 19610 23136 19612
rect 23160 19610 23216 19612
rect 23240 19610 23296 19612
rect 22920 19558 22922 19610
rect 22922 19558 22974 19610
rect 22974 19558 22976 19610
rect 23000 19558 23038 19610
rect 23038 19558 23050 19610
rect 23050 19558 23056 19610
rect 23080 19558 23102 19610
rect 23102 19558 23114 19610
rect 23114 19558 23136 19610
rect 23160 19558 23166 19610
rect 23166 19558 23178 19610
rect 23178 19558 23216 19610
rect 23240 19558 23242 19610
rect 23242 19558 23294 19610
rect 23294 19558 23296 19610
rect 22920 19556 22976 19558
rect 23000 19556 23056 19558
rect 23080 19556 23136 19558
rect 23160 19556 23216 19558
rect 23240 19556 23296 19558
rect 28180 27770 28236 27772
rect 28260 27770 28316 27772
rect 28340 27770 28396 27772
rect 28420 27770 28476 27772
rect 28500 27770 28556 27772
rect 28180 27718 28182 27770
rect 28182 27718 28234 27770
rect 28234 27718 28236 27770
rect 28260 27718 28298 27770
rect 28298 27718 28310 27770
rect 28310 27718 28316 27770
rect 28340 27718 28362 27770
rect 28362 27718 28374 27770
rect 28374 27718 28396 27770
rect 28420 27718 28426 27770
rect 28426 27718 28438 27770
rect 28438 27718 28476 27770
rect 28500 27718 28502 27770
rect 28502 27718 28554 27770
rect 28554 27718 28556 27770
rect 28180 27716 28236 27718
rect 28260 27716 28316 27718
rect 28340 27716 28396 27718
rect 28420 27716 28476 27718
rect 28500 27716 28556 27718
rect 24858 21564 24860 21584
rect 24860 21564 24912 21584
rect 24912 21564 24914 21584
rect 24858 21528 24914 21564
rect 22180 17978 22236 17980
rect 22260 17978 22316 17980
rect 22340 17978 22396 17980
rect 22420 17978 22476 17980
rect 22500 17978 22556 17980
rect 22180 17926 22182 17978
rect 22182 17926 22234 17978
rect 22234 17926 22236 17978
rect 22260 17926 22298 17978
rect 22298 17926 22310 17978
rect 22310 17926 22316 17978
rect 22340 17926 22362 17978
rect 22362 17926 22374 17978
rect 22374 17926 22396 17978
rect 22420 17926 22426 17978
rect 22426 17926 22438 17978
rect 22438 17926 22476 17978
rect 22500 17926 22502 17978
rect 22502 17926 22554 17978
rect 22554 17926 22556 17978
rect 22180 17924 22236 17926
rect 22260 17924 22316 17926
rect 22340 17924 22396 17926
rect 22420 17924 22476 17926
rect 22500 17924 22556 17926
rect 22180 16890 22236 16892
rect 22260 16890 22316 16892
rect 22340 16890 22396 16892
rect 22420 16890 22476 16892
rect 22500 16890 22556 16892
rect 22180 16838 22182 16890
rect 22182 16838 22234 16890
rect 22234 16838 22236 16890
rect 22260 16838 22298 16890
rect 22298 16838 22310 16890
rect 22310 16838 22316 16890
rect 22340 16838 22362 16890
rect 22362 16838 22374 16890
rect 22374 16838 22396 16890
rect 22420 16838 22426 16890
rect 22426 16838 22438 16890
rect 22438 16838 22476 16890
rect 22500 16838 22502 16890
rect 22502 16838 22554 16890
rect 22554 16838 22556 16890
rect 22180 16836 22236 16838
rect 22260 16836 22316 16838
rect 22340 16836 22396 16838
rect 22420 16836 22476 16838
rect 22500 16836 22556 16838
rect 21362 15988 21364 16008
rect 21364 15988 21416 16008
rect 21416 15988 21418 16008
rect 21362 15952 21418 15988
rect 16920 5466 16976 5468
rect 17000 5466 17056 5468
rect 17080 5466 17136 5468
rect 17160 5466 17216 5468
rect 17240 5466 17296 5468
rect 16920 5414 16922 5466
rect 16922 5414 16974 5466
rect 16974 5414 16976 5466
rect 17000 5414 17038 5466
rect 17038 5414 17050 5466
rect 17050 5414 17056 5466
rect 17080 5414 17102 5466
rect 17102 5414 17114 5466
rect 17114 5414 17136 5466
rect 17160 5414 17166 5466
rect 17166 5414 17178 5466
rect 17178 5414 17216 5466
rect 17240 5414 17242 5466
rect 17242 5414 17294 5466
rect 17294 5414 17296 5466
rect 16920 5412 16976 5414
rect 17000 5412 17056 5414
rect 17080 5412 17136 5414
rect 17160 5412 17216 5414
rect 17240 5412 17296 5414
rect 20442 12688 20498 12744
rect 21638 11772 21640 11792
rect 21640 11772 21692 11792
rect 21692 11772 21694 11792
rect 21638 11736 21694 11772
rect 16180 4922 16236 4924
rect 16260 4922 16316 4924
rect 16340 4922 16396 4924
rect 16420 4922 16476 4924
rect 16500 4922 16556 4924
rect 16180 4870 16182 4922
rect 16182 4870 16234 4922
rect 16234 4870 16236 4922
rect 16260 4870 16298 4922
rect 16298 4870 16310 4922
rect 16310 4870 16316 4922
rect 16340 4870 16362 4922
rect 16362 4870 16374 4922
rect 16374 4870 16396 4922
rect 16420 4870 16426 4922
rect 16426 4870 16438 4922
rect 16438 4870 16476 4922
rect 16500 4870 16502 4922
rect 16502 4870 16554 4922
rect 16554 4870 16556 4922
rect 16180 4868 16236 4870
rect 16260 4868 16316 4870
rect 16340 4868 16396 4870
rect 16420 4868 16476 4870
rect 16500 4868 16556 4870
rect 22180 15802 22236 15804
rect 22260 15802 22316 15804
rect 22340 15802 22396 15804
rect 22420 15802 22476 15804
rect 22500 15802 22556 15804
rect 22180 15750 22182 15802
rect 22182 15750 22234 15802
rect 22234 15750 22236 15802
rect 22260 15750 22298 15802
rect 22298 15750 22310 15802
rect 22310 15750 22316 15802
rect 22340 15750 22362 15802
rect 22362 15750 22374 15802
rect 22374 15750 22396 15802
rect 22420 15750 22426 15802
rect 22426 15750 22438 15802
rect 22438 15750 22476 15802
rect 22500 15750 22502 15802
rect 22502 15750 22554 15802
rect 22554 15750 22556 15802
rect 22180 15748 22236 15750
rect 22260 15748 22316 15750
rect 22340 15748 22396 15750
rect 22420 15748 22476 15750
rect 22500 15748 22556 15750
rect 22180 14714 22236 14716
rect 22260 14714 22316 14716
rect 22340 14714 22396 14716
rect 22420 14714 22476 14716
rect 22500 14714 22556 14716
rect 22180 14662 22182 14714
rect 22182 14662 22234 14714
rect 22234 14662 22236 14714
rect 22260 14662 22298 14714
rect 22298 14662 22310 14714
rect 22310 14662 22316 14714
rect 22340 14662 22362 14714
rect 22362 14662 22374 14714
rect 22374 14662 22396 14714
rect 22420 14662 22426 14714
rect 22426 14662 22438 14714
rect 22438 14662 22476 14714
rect 22500 14662 22502 14714
rect 22502 14662 22554 14714
rect 22554 14662 22556 14714
rect 22180 14660 22236 14662
rect 22260 14660 22316 14662
rect 22340 14660 22396 14662
rect 22420 14660 22476 14662
rect 22500 14660 22556 14662
rect 22180 13626 22236 13628
rect 22260 13626 22316 13628
rect 22340 13626 22396 13628
rect 22420 13626 22476 13628
rect 22500 13626 22556 13628
rect 22180 13574 22182 13626
rect 22182 13574 22234 13626
rect 22234 13574 22236 13626
rect 22260 13574 22298 13626
rect 22298 13574 22310 13626
rect 22310 13574 22316 13626
rect 22340 13574 22362 13626
rect 22362 13574 22374 13626
rect 22374 13574 22396 13626
rect 22420 13574 22426 13626
rect 22426 13574 22438 13626
rect 22438 13574 22476 13626
rect 22500 13574 22502 13626
rect 22502 13574 22554 13626
rect 22554 13574 22556 13626
rect 22180 13572 22236 13574
rect 22260 13572 22316 13574
rect 22340 13572 22396 13574
rect 22420 13572 22476 13574
rect 22500 13572 22556 13574
rect 22180 12538 22236 12540
rect 22260 12538 22316 12540
rect 22340 12538 22396 12540
rect 22420 12538 22476 12540
rect 22500 12538 22556 12540
rect 22180 12486 22182 12538
rect 22182 12486 22234 12538
rect 22234 12486 22236 12538
rect 22260 12486 22298 12538
rect 22298 12486 22310 12538
rect 22310 12486 22316 12538
rect 22340 12486 22362 12538
rect 22362 12486 22374 12538
rect 22374 12486 22396 12538
rect 22420 12486 22426 12538
rect 22426 12486 22438 12538
rect 22438 12486 22476 12538
rect 22500 12486 22502 12538
rect 22502 12486 22554 12538
rect 22554 12486 22556 12538
rect 22180 12484 22236 12486
rect 22260 12484 22316 12486
rect 22340 12484 22396 12486
rect 22420 12484 22476 12486
rect 22500 12484 22556 12486
rect 22180 11450 22236 11452
rect 22260 11450 22316 11452
rect 22340 11450 22396 11452
rect 22420 11450 22476 11452
rect 22500 11450 22556 11452
rect 22180 11398 22182 11450
rect 22182 11398 22234 11450
rect 22234 11398 22236 11450
rect 22260 11398 22298 11450
rect 22298 11398 22310 11450
rect 22310 11398 22316 11450
rect 22340 11398 22362 11450
rect 22362 11398 22374 11450
rect 22374 11398 22396 11450
rect 22420 11398 22426 11450
rect 22426 11398 22438 11450
rect 22438 11398 22476 11450
rect 22500 11398 22502 11450
rect 22502 11398 22554 11450
rect 22554 11398 22556 11450
rect 22180 11396 22236 11398
rect 22260 11396 22316 11398
rect 22340 11396 22396 11398
rect 22420 11396 22476 11398
rect 22500 11396 22556 11398
rect 22180 10362 22236 10364
rect 22260 10362 22316 10364
rect 22340 10362 22396 10364
rect 22420 10362 22476 10364
rect 22500 10362 22556 10364
rect 22180 10310 22182 10362
rect 22182 10310 22234 10362
rect 22234 10310 22236 10362
rect 22260 10310 22298 10362
rect 22298 10310 22310 10362
rect 22310 10310 22316 10362
rect 22340 10310 22362 10362
rect 22362 10310 22374 10362
rect 22374 10310 22396 10362
rect 22420 10310 22426 10362
rect 22426 10310 22438 10362
rect 22438 10310 22476 10362
rect 22500 10310 22502 10362
rect 22502 10310 22554 10362
rect 22554 10310 22556 10362
rect 22180 10308 22236 10310
rect 22260 10308 22316 10310
rect 22340 10308 22396 10310
rect 22420 10308 22476 10310
rect 22500 10308 22556 10310
rect 22180 9274 22236 9276
rect 22260 9274 22316 9276
rect 22340 9274 22396 9276
rect 22420 9274 22476 9276
rect 22500 9274 22556 9276
rect 22180 9222 22182 9274
rect 22182 9222 22234 9274
rect 22234 9222 22236 9274
rect 22260 9222 22298 9274
rect 22298 9222 22310 9274
rect 22310 9222 22316 9274
rect 22340 9222 22362 9274
rect 22362 9222 22374 9274
rect 22374 9222 22396 9274
rect 22420 9222 22426 9274
rect 22426 9222 22438 9274
rect 22438 9222 22476 9274
rect 22500 9222 22502 9274
rect 22502 9222 22554 9274
rect 22554 9222 22556 9274
rect 22180 9220 22236 9222
rect 22260 9220 22316 9222
rect 22340 9220 22396 9222
rect 22420 9220 22476 9222
rect 22500 9220 22556 9222
rect 22920 18522 22976 18524
rect 23000 18522 23056 18524
rect 23080 18522 23136 18524
rect 23160 18522 23216 18524
rect 23240 18522 23296 18524
rect 22920 18470 22922 18522
rect 22922 18470 22974 18522
rect 22974 18470 22976 18522
rect 23000 18470 23038 18522
rect 23038 18470 23050 18522
rect 23050 18470 23056 18522
rect 23080 18470 23102 18522
rect 23102 18470 23114 18522
rect 23114 18470 23136 18522
rect 23160 18470 23166 18522
rect 23166 18470 23178 18522
rect 23178 18470 23216 18522
rect 23240 18470 23242 18522
rect 23242 18470 23294 18522
rect 23294 18470 23296 18522
rect 22920 18468 22976 18470
rect 23000 18468 23056 18470
rect 23080 18468 23136 18470
rect 23160 18468 23216 18470
rect 23240 18468 23296 18470
rect 22920 17434 22976 17436
rect 23000 17434 23056 17436
rect 23080 17434 23136 17436
rect 23160 17434 23216 17436
rect 23240 17434 23296 17436
rect 22920 17382 22922 17434
rect 22922 17382 22974 17434
rect 22974 17382 22976 17434
rect 23000 17382 23038 17434
rect 23038 17382 23050 17434
rect 23050 17382 23056 17434
rect 23080 17382 23102 17434
rect 23102 17382 23114 17434
rect 23114 17382 23136 17434
rect 23160 17382 23166 17434
rect 23166 17382 23178 17434
rect 23178 17382 23216 17434
rect 23240 17382 23242 17434
rect 23242 17382 23294 17434
rect 23294 17382 23296 17434
rect 22920 17380 22976 17382
rect 23000 17380 23056 17382
rect 23080 17380 23136 17382
rect 23160 17380 23216 17382
rect 23240 17380 23296 17382
rect 22920 16346 22976 16348
rect 23000 16346 23056 16348
rect 23080 16346 23136 16348
rect 23160 16346 23216 16348
rect 23240 16346 23296 16348
rect 22920 16294 22922 16346
rect 22922 16294 22974 16346
rect 22974 16294 22976 16346
rect 23000 16294 23038 16346
rect 23038 16294 23050 16346
rect 23050 16294 23056 16346
rect 23080 16294 23102 16346
rect 23102 16294 23114 16346
rect 23114 16294 23136 16346
rect 23160 16294 23166 16346
rect 23166 16294 23178 16346
rect 23178 16294 23216 16346
rect 23240 16294 23242 16346
rect 23242 16294 23294 16346
rect 23294 16294 23296 16346
rect 22920 16292 22976 16294
rect 23000 16292 23056 16294
rect 23080 16292 23136 16294
rect 23160 16292 23216 16294
rect 23240 16292 23296 16294
rect 22926 15952 22982 16008
rect 22920 15258 22976 15260
rect 23000 15258 23056 15260
rect 23080 15258 23136 15260
rect 23160 15258 23216 15260
rect 23240 15258 23296 15260
rect 22920 15206 22922 15258
rect 22922 15206 22974 15258
rect 22974 15206 22976 15258
rect 23000 15206 23038 15258
rect 23038 15206 23050 15258
rect 23050 15206 23056 15258
rect 23080 15206 23102 15258
rect 23102 15206 23114 15258
rect 23114 15206 23136 15258
rect 23160 15206 23166 15258
rect 23166 15206 23178 15258
rect 23178 15206 23216 15258
rect 23240 15206 23242 15258
rect 23242 15206 23294 15258
rect 23294 15206 23296 15258
rect 22920 15204 22976 15206
rect 23000 15204 23056 15206
rect 23080 15204 23136 15206
rect 23160 15204 23216 15206
rect 23240 15204 23296 15206
rect 22920 14170 22976 14172
rect 23000 14170 23056 14172
rect 23080 14170 23136 14172
rect 23160 14170 23216 14172
rect 23240 14170 23296 14172
rect 22920 14118 22922 14170
rect 22922 14118 22974 14170
rect 22974 14118 22976 14170
rect 23000 14118 23038 14170
rect 23038 14118 23050 14170
rect 23050 14118 23056 14170
rect 23080 14118 23102 14170
rect 23102 14118 23114 14170
rect 23114 14118 23136 14170
rect 23160 14118 23166 14170
rect 23166 14118 23178 14170
rect 23178 14118 23216 14170
rect 23240 14118 23242 14170
rect 23242 14118 23294 14170
rect 23294 14118 23296 14170
rect 22920 14116 22976 14118
rect 23000 14116 23056 14118
rect 23080 14116 23136 14118
rect 23160 14116 23216 14118
rect 23240 14116 23296 14118
rect 22920 13082 22976 13084
rect 23000 13082 23056 13084
rect 23080 13082 23136 13084
rect 23160 13082 23216 13084
rect 23240 13082 23296 13084
rect 22920 13030 22922 13082
rect 22922 13030 22974 13082
rect 22974 13030 22976 13082
rect 23000 13030 23038 13082
rect 23038 13030 23050 13082
rect 23050 13030 23056 13082
rect 23080 13030 23102 13082
rect 23102 13030 23114 13082
rect 23114 13030 23136 13082
rect 23160 13030 23166 13082
rect 23166 13030 23178 13082
rect 23178 13030 23216 13082
rect 23240 13030 23242 13082
rect 23242 13030 23294 13082
rect 23294 13030 23296 13082
rect 22920 13028 22976 13030
rect 23000 13028 23056 13030
rect 23080 13028 23136 13030
rect 23160 13028 23216 13030
rect 23240 13028 23296 13030
rect 22920 11994 22976 11996
rect 23000 11994 23056 11996
rect 23080 11994 23136 11996
rect 23160 11994 23216 11996
rect 23240 11994 23296 11996
rect 22920 11942 22922 11994
rect 22922 11942 22974 11994
rect 22974 11942 22976 11994
rect 23000 11942 23038 11994
rect 23038 11942 23050 11994
rect 23050 11942 23056 11994
rect 23080 11942 23102 11994
rect 23102 11942 23114 11994
rect 23114 11942 23136 11994
rect 23160 11942 23166 11994
rect 23166 11942 23178 11994
rect 23178 11942 23216 11994
rect 23240 11942 23242 11994
rect 23242 11942 23294 11994
rect 23294 11942 23296 11994
rect 22920 11940 22976 11942
rect 23000 11940 23056 11942
rect 23080 11940 23136 11942
rect 23160 11940 23216 11942
rect 23240 11940 23296 11942
rect 22920 10906 22976 10908
rect 23000 10906 23056 10908
rect 23080 10906 23136 10908
rect 23160 10906 23216 10908
rect 23240 10906 23296 10908
rect 22920 10854 22922 10906
rect 22922 10854 22974 10906
rect 22974 10854 22976 10906
rect 23000 10854 23038 10906
rect 23038 10854 23050 10906
rect 23050 10854 23056 10906
rect 23080 10854 23102 10906
rect 23102 10854 23114 10906
rect 23114 10854 23136 10906
rect 23160 10854 23166 10906
rect 23166 10854 23178 10906
rect 23178 10854 23216 10906
rect 23240 10854 23242 10906
rect 23242 10854 23294 10906
rect 23294 10854 23296 10906
rect 22920 10852 22976 10854
rect 23000 10852 23056 10854
rect 23080 10852 23136 10854
rect 23160 10852 23216 10854
rect 23240 10852 23296 10854
rect 22920 9818 22976 9820
rect 23000 9818 23056 9820
rect 23080 9818 23136 9820
rect 23160 9818 23216 9820
rect 23240 9818 23296 9820
rect 22920 9766 22922 9818
rect 22922 9766 22974 9818
rect 22974 9766 22976 9818
rect 23000 9766 23038 9818
rect 23038 9766 23050 9818
rect 23050 9766 23056 9818
rect 23080 9766 23102 9818
rect 23102 9766 23114 9818
rect 23114 9766 23136 9818
rect 23160 9766 23166 9818
rect 23166 9766 23178 9818
rect 23178 9766 23216 9818
rect 23240 9766 23242 9818
rect 23242 9766 23294 9818
rect 23294 9766 23296 9818
rect 22920 9764 22976 9766
rect 23000 9764 23056 9766
rect 23080 9764 23136 9766
rect 23160 9764 23216 9766
rect 23240 9764 23296 9766
rect 28920 27226 28976 27228
rect 29000 27226 29056 27228
rect 29080 27226 29136 27228
rect 29160 27226 29216 27228
rect 29240 27226 29296 27228
rect 28920 27174 28922 27226
rect 28922 27174 28974 27226
rect 28974 27174 28976 27226
rect 29000 27174 29038 27226
rect 29038 27174 29050 27226
rect 29050 27174 29056 27226
rect 29080 27174 29102 27226
rect 29102 27174 29114 27226
rect 29114 27174 29136 27226
rect 29160 27174 29166 27226
rect 29166 27174 29178 27226
rect 29178 27174 29216 27226
rect 29240 27174 29242 27226
rect 29242 27174 29294 27226
rect 29294 27174 29296 27226
rect 28920 27172 28976 27174
rect 29000 27172 29056 27174
rect 29080 27172 29136 27174
rect 29160 27172 29216 27174
rect 29240 27172 29296 27174
rect 23846 15952 23902 16008
rect 28180 26682 28236 26684
rect 28260 26682 28316 26684
rect 28340 26682 28396 26684
rect 28420 26682 28476 26684
rect 28500 26682 28556 26684
rect 28180 26630 28182 26682
rect 28182 26630 28234 26682
rect 28234 26630 28236 26682
rect 28260 26630 28298 26682
rect 28298 26630 28310 26682
rect 28310 26630 28316 26682
rect 28340 26630 28362 26682
rect 28362 26630 28374 26682
rect 28374 26630 28396 26682
rect 28420 26630 28426 26682
rect 28426 26630 28438 26682
rect 28438 26630 28476 26682
rect 28500 26630 28502 26682
rect 28502 26630 28554 26682
rect 28554 26630 28556 26682
rect 28180 26628 28236 26630
rect 28260 26628 28316 26630
rect 28340 26628 28396 26630
rect 28420 26628 28476 26630
rect 28500 26628 28556 26630
rect 28920 26138 28976 26140
rect 29000 26138 29056 26140
rect 29080 26138 29136 26140
rect 29160 26138 29216 26140
rect 29240 26138 29296 26140
rect 28920 26086 28922 26138
rect 28922 26086 28974 26138
rect 28974 26086 28976 26138
rect 29000 26086 29038 26138
rect 29038 26086 29050 26138
rect 29050 26086 29056 26138
rect 29080 26086 29102 26138
rect 29102 26086 29114 26138
rect 29114 26086 29136 26138
rect 29160 26086 29166 26138
rect 29166 26086 29178 26138
rect 29178 26086 29216 26138
rect 29240 26086 29242 26138
rect 29242 26086 29294 26138
rect 29294 26086 29296 26138
rect 28920 26084 28976 26086
rect 29000 26084 29056 26086
rect 29080 26084 29136 26086
rect 29160 26084 29216 26086
rect 29240 26084 29296 26086
rect 28180 25594 28236 25596
rect 28260 25594 28316 25596
rect 28340 25594 28396 25596
rect 28420 25594 28476 25596
rect 28500 25594 28556 25596
rect 28180 25542 28182 25594
rect 28182 25542 28234 25594
rect 28234 25542 28236 25594
rect 28260 25542 28298 25594
rect 28298 25542 28310 25594
rect 28310 25542 28316 25594
rect 28340 25542 28362 25594
rect 28362 25542 28374 25594
rect 28374 25542 28396 25594
rect 28420 25542 28426 25594
rect 28426 25542 28438 25594
rect 28438 25542 28476 25594
rect 28500 25542 28502 25594
rect 28502 25542 28554 25594
rect 28554 25542 28556 25594
rect 28180 25540 28236 25542
rect 28260 25540 28316 25542
rect 28340 25540 28396 25542
rect 28420 25540 28476 25542
rect 28500 25540 28556 25542
rect 28920 25050 28976 25052
rect 29000 25050 29056 25052
rect 29080 25050 29136 25052
rect 29160 25050 29216 25052
rect 29240 25050 29296 25052
rect 28920 24998 28922 25050
rect 28922 24998 28974 25050
rect 28974 24998 28976 25050
rect 29000 24998 29038 25050
rect 29038 24998 29050 25050
rect 29050 24998 29056 25050
rect 29080 24998 29102 25050
rect 29102 24998 29114 25050
rect 29114 24998 29136 25050
rect 29160 24998 29166 25050
rect 29166 24998 29178 25050
rect 29178 24998 29216 25050
rect 29240 24998 29242 25050
rect 29242 24998 29294 25050
rect 29294 24998 29296 25050
rect 28920 24996 28976 24998
rect 29000 24996 29056 24998
rect 29080 24996 29136 24998
rect 29160 24996 29216 24998
rect 29240 24996 29296 24998
rect 28180 24506 28236 24508
rect 28260 24506 28316 24508
rect 28340 24506 28396 24508
rect 28420 24506 28476 24508
rect 28500 24506 28556 24508
rect 28180 24454 28182 24506
rect 28182 24454 28234 24506
rect 28234 24454 28236 24506
rect 28260 24454 28298 24506
rect 28298 24454 28310 24506
rect 28310 24454 28316 24506
rect 28340 24454 28362 24506
rect 28362 24454 28374 24506
rect 28374 24454 28396 24506
rect 28420 24454 28426 24506
rect 28426 24454 28438 24506
rect 28438 24454 28476 24506
rect 28500 24454 28502 24506
rect 28502 24454 28554 24506
rect 28554 24454 28556 24506
rect 28180 24452 28236 24454
rect 28260 24452 28316 24454
rect 28340 24452 28396 24454
rect 28420 24452 28476 24454
rect 28500 24452 28556 24454
rect 28920 23962 28976 23964
rect 29000 23962 29056 23964
rect 29080 23962 29136 23964
rect 29160 23962 29216 23964
rect 29240 23962 29296 23964
rect 28920 23910 28922 23962
rect 28922 23910 28974 23962
rect 28974 23910 28976 23962
rect 29000 23910 29038 23962
rect 29038 23910 29050 23962
rect 29050 23910 29056 23962
rect 29080 23910 29102 23962
rect 29102 23910 29114 23962
rect 29114 23910 29136 23962
rect 29160 23910 29166 23962
rect 29166 23910 29178 23962
rect 29178 23910 29216 23962
rect 29240 23910 29242 23962
rect 29242 23910 29294 23962
rect 29294 23910 29296 23962
rect 28920 23908 28976 23910
rect 29000 23908 29056 23910
rect 29080 23908 29136 23910
rect 29160 23908 29216 23910
rect 29240 23908 29296 23910
rect 28180 23418 28236 23420
rect 28260 23418 28316 23420
rect 28340 23418 28396 23420
rect 28420 23418 28476 23420
rect 28500 23418 28556 23420
rect 28180 23366 28182 23418
rect 28182 23366 28234 23418
rect 28234 23366 28236 23418
rect 28260 23366 28298 23418
rect 28298 23366 28310 23418
rect 28310 23366 28316 23418
rect 28340 23366 28362 23418
rect 28362 23366 28374 23418
rect 28374 23366 28396 23418
rect 28420 23366 28426 23418
rect 28426 23366 28438 23418
rect 28438 23366 28476 23418
rect 28500 23366 28502 23418
rect 28502 23366 28554 23418
rect 28554 23366 28556 23418
rect 28180 23364 28236 23366
rect 28260 23364 28316 23366
rect 28340 23364 28396 23366
rect 28420 23364 28476 23366
rect 28500 23364 28556 23366
rect 28180 22330 28236 22332
rect 28260 22330 28316 22332
rect 28340 22330 28396 22332
rect 28420 22330 28476 22332
rect 28500 22330 28556 22332
rect 28180 22278 28182 22330
rect 28182 22278 28234 22330
rect 28234 22278 28236 22330
rect 28260 22278 28298 22330
rect 28298 22278 28310 22330
rect 28310 22278 28316 22330
rect 28340 22278 28362 22330
rect 28362 22278 28374 22330
rect 28374 22278 28396 22330
rect 28420 22278 28426 22330
rect 28426 22278 28438 22330
rect 28438 22278 28476 22330
rect 28500 22278 28502 22330
rect 28502 22278 28554 22330
rect 28554 22278 28556 22330
rect 28180 22276 28236 22278
rect 28260 22276 28316 22278
rect 28340 22276 28396 22278
rect 28420 22276 28476 22278
rect 28500 22276 28556 22278
rect 28180 21242 28236 21244
rect 28260 21242 28316 21244
rect 28340 21242 28396 21244
rect 28420 21242 28476 21244
rect 28500 21242 28556 21244
rect 28180 21190 28182 21242
rect 28182 21190 28234 21242
rect 28234 21190 28236 21242
rect 28260 21190 28298 21242
rect 28298 21190 28310 21242
rect 28310 21190 28316 21242
rect 28340 21190 28362 21242
rect 28362 21190 28374 21242
rect 28374 21190 28396 21242
rect 28420 21190 28426 21242
rect 28426 21190 28438 21242
rect 28438 21190 28476 21242
rect 28500 21190 28502 21242
rect 28502 21190 28554 21242
rect 28554 21190 28556 21242
rect 28180 21188 28236 21190
rect 28260 21188 28316 21190
rect 28340 21188 28396 21190
rect 28420 21188 28476 21190
rect 28500 21188 28556 21190
rect 28180 20154 28236 20156
rect 28260 20154 28316 20156
rect 28340 20154 28396 20156
rect 28420 20154 28476 20156
rect 28500 20154 28556 20156
rect 28180 20102 28182 20154
rect 28182 20102 28234 20154
rect 28234 20102 28236 20154
rect 28260 20102 28298 20154
rect 28298 20102 28310 20154
rect 28310 20102 28316 20154
rect 28340 20102 28362 20154
rect 28362 20102 28374 20154
rect 28374 20102 28396 20154
rect 28420 20102 28426 20154
rect 28426 20102 28438 20154
rect 28438 20102 28476 20154
rect 28500 20102 28502 20154
rect 28502 20102 28554 20154
rect 28554 20102 28556 20154
rect 28180 20100 28236 20102
rect 28260 20100 28316 20102
rect 28340 20100 28396 20102
rect 28420 20100 28476 20102
rect 28500 20100 28556 20102
rect 28920 22874 28976 22876
rect 29000 22874 29056 22876
rect 29080 22874 29136 22876
rect 29160 22874 29216 22876
rect 29240 22874 29296 22876
rect 28920 22822 28922 22874
rect 28922 22822 28974 22874
rect 28974 22822 28976 22874
rect 29000 22822 29038 22874
rect 29038 22822 29050 22874
rect 29050 22822 29056 22874
rect 29080 22822 29102 22874
rect 29102 22822 29114 22874
rect 29114 22822 29136 22874
rect 29160 22822 29166 22874
rect 29166 22822 29178 22874
rect 29178 22822 29216 22874
rect 29240 22822 29242 22874
rect 29242 22822 29294 22874
rect 29294 22822 29296 22874
rect 28920 22820 28976 22822
rect 29000 22820 29056 22822
rect 29080 22820 29136 22822
rect 29160 22820 29216 22822
rect 29240 22820 29296 22822
rect 28920 21786 28976 21788
rect 29000 21786 29056 21788
rect 29080 21786 29136 21788
rect 29160 21786 29216 21788
rect 29240 21786 29296 21788
rect 28920 21734 28922 21786
rect 28922 21734 28974 21786
rect 28974 21734 28976 21786
rect 29000 21734 29038 21786
rect 29038 21734 29050 21786
rect 29050 21734 29056 21786
rect 29080 21734 29102 21786
rect 29102 21734 29114 21786
rect 29114 21734 29136 21786
rect 29160 21734 29166 21786
rect 29166 21734 29178 21786
rect 29178 21734 29216 21786
rect 29240 21734 29242 21786
rect 29242 21734 29294 21786
rect 29294 21734 29296 21786
rect 28920 21732 28976 21734
rect 29000 21732 29056 21734
rect 29080 21732 29136 21734
rect 29160 21732 29216 21734
rect 29240 21732 29296 21734
rect 28920 20698 28976 20700
rect 29000 20698 29056 20700
rect 29080 20698 29136 20700
rect 29160 20698 29216 20700
rect 29240 20698 29296 20700
rect 28920 20646 28922 20698
rect 28922 20646 28974 20698
rect 28974 20646 28976 20698
rect 29000 20646 29038 20698
rect 29038 20646 29050 20698
rect 29050 20646 29056 20698
rect 29080 20646 29102 20698
rect 29102 20646 29114 20698
rect 29114 20646 29136 20698
rect 29160 20646 29166 20698
rect 29166 20646 29178 20698
rect 29178 20646 29216 20698
rect 29240 20646 29242 20698
rect 29242 20646 29294 20698
rect 29294 20646 29296 20698
rect 28920 20644 28976 20646
rect 29000 20644 29056 20646
rect 29080 20644 29136 20646
rect 29160 20644 29216 20646
rect 29240 20644 29296 20646
rect 31482 25880 31538 25936
rect 31114 24656 31170 24712
rect 28920 19610 28976 19612
rect 29000 19610 29056 19612
rect 29080 19610 29136 19612
rect 29160 19610 29216 19612
rect 29240 19610 29296 19612
rect 28920 19558 28922 19610
rect 28922 19558 28974 19610
rect 28974 19558 28976 19610
rect 29000 19558 29038 19610
rect 29038 19558 29050 19610
rect 29050 19558 29056 19610
rect 29080 19558 29102 19610
rect 29102 19558 29114 19610
rect 29114 19558 29136 19610
rect 29160 19558 29166 19610
rect 29166 19558 29178 19610
rect 29178 19558 29216 19610
rect 29240 19558 29242 19610
rect 29242 19558 29294 19610
rect 29294 19558 29296 19610
rect 28920 19556 28976 19558
rect 29000 19556 29056 19558
rect 29080 19556 29136 19558
rect 29160 19556 29216 19558
rect 29240 19556 29296 19558
rect 28180 19066 28236 19068
rect 28260 19066 28316 19068
rect 28340 19066 28396 19068
rect 28420 19066 28476 19068
rect 28500 19066 28556 19068
rect 28180 19014 28182 19066
rect 28182 19014 28234 19066
rect 28234 19014 28236 19066
rect 28260 19014 28298 19066
rect 28298 19014 28310 19066
rect 28310 19014 28316 19066
rect 28340 19014 28362 19066
rect 28362 19014 28374 19066
rect 28374 19014 28396 19066
rect 28420 19014 28426 19066
rect 28426 19014 28438 19066
rect 28438 19014 28476 19066
rect 28500 19014 28502 19066
rect 28502 19014 28554 19066
rect 28554 19014 28556 19066
rect 28180 19012 28236 19014
rect 28260 19012 28316 19014
rect 28340 19012 28396 19014
rect 28420 19012 28476 19014
rect 28500 19012 28556 19014
rect 28920 18522 28976 18524
rect 29000 18522 29056 18524
rect 29080 18522 29136 18524
rect 29160 18522 29216 18524
rect 29240 18522 29296 18524
rect 28920 18470 28922 18522
rect 28922 18470 28974 18522
rect 28974 18470 28976 18522
rect 29000 18470 29038 18522
rect 29038 18470 29050 18522
rect 29050 18470 29056 18522
rect 29080 18470 29102 18522
rect 29102 18470 29114 18522
rect 29114 18470 29136 18522
rect 29160 18470 29166 18522
rect 29166 18470 29178 18522
rect 29178 18470 29216 18522
rect 29240 18470 29242 18522
rect 29242 18470 29294 18522
rect 29294 18470 29296 18522
rect 28920 18468 28976 18470
rect 29000 18468 29056 18470
rect 29080 18468 29136 18470
rect 29160 18468 29216 18470
rect 29240 18468 29296 18470
rect 28180 17978 28236 17980
rect 28260 17978 28316 17980
rect 28340 17978 28396 17980
rect 28420 17978 28476 17980
rect 28500 17978 28556 17980
rect 28180 17926 28182 17978
rect 28182 17926 28234 17978
rect 28234 17926 28236 17978
rect 28260 17926 28298 17978
rect 28298 17926 28310 17978
rect 28310 17926 28316 17978
rect 28340 17926 28362 17978
rect 28362 17926 28374 17978
rect 28374 17926 28396 17978
rect 28420 17926 28426 17978
rect 28426 17926 28438 17978
rect 28438 17926 28476 17978
rect 28500 17926 28502 17978
rect 28502 17926 28554 17978
rect 28554 17926 28556 17978
rect 28180 17924 28236 17926
rect 28260 17924 28316 17926
rect 28340 17924 28396 17926
rect 28420 17924 28476 17926
rect 28500 17924 28556 17926
rect 28920 17434 28976 17436
rect 29000 17434 29056 17436
rect 29080 17434 29136 17436
rect 29160 17434 29216 17436
rect 29240 17434 29296 17436
rect 28920 17382 28922 17434
rect 28922 17382 28974 17434
rect 28974 17382 28976 17434
rect 29000 17382 29038 17434
rect 29038 17382 29050 17434
rect 29050 17382 29056 17434
rect 29080 17382 29102 17434
rect 29102 17382 29114 17434
rect 29114 17382 29136 17434
rect 29160 17382 29166 17434
rect 29166 17382 29178 17434
rect 29178 17382 29216 17434
rect 29240 17382 29242 17434
rect 29242 17382 29294 17434
rect 29294 17382 29296 17434
rect 28920 17380 28976 17382
rect 29000 17380 29056 17382
rect 29080 17380 29136 17382
rect 29160 17380 29216 17382
rect 29240 17380 29296 17382
rect 28180 16890 28236 16892
rect 28260 16890 28316 16892
rect 28340 16890 28396 16892
rect 28420 16890 28476 16892
rect 28500 16890 28556 16892
rect 28180 16838 28182 16890
rect 28182 16838 28234 16890
rect 28234 16838 28236 16890
rect 28260 16838 28298 16890
rect 28298 16838 28310 16890
rect 28310 16838 28316 16890
rect 28340 16838 28362 16890
rect 28362 16838 28374 16890
rect 28374 16838 28396 16890
rect 28420 16838 28426 16890
rect 28426 16838 28438 16890
rect 28438 16838 28476 16890
rect 28500 16838 28502 16890
rect 28502 16838 28554 16890
rect 28554 16838 28556 16890
rect 28180 16836 28236 16838
rect 28260 16836 28316 16838
rect 28340 16836 28396 16838
rect 28420 16836 28476 16838
rect 28500 16836 28556 16838
rect 25410 11736 25466 11792
rect 22180 8186 22236 8188
rect 22260 8186 22316 8188
rect 22340 8186 22396 8188
rect 22420 8186 22476 8188
rect 22500 8186 22556 8188
rect 22180 8134 22182 8186
rect 22182 8134 22234 8186
rect 22234 8134 22236 8186
rect 22260 8134 22298 8186
rect 22298 8134 22310 8186
rect 22310 8134 22316 8186
rect 22340 8134 22362 8186
rect 22362 8134 22374 8186
rect 22374 8134 22396 8186
rect 22420 8134 22426 8186
rect 22426 8134 22438 8186
rect 22438 8134 22476 8186
rect 22500 8134 22502 8186
rect 22502 8134 22554 8186
rect 22554 8134 22556 8186
rect 22180 8132 22236 8134
rect 22260 8132 22316 8134
rect 22340 8132 22396 8134
rect 22420 8132 22476 8134
rect 22500 8132 22556 8134
rect 22180 7098 22236 7100
rect 22260 7098 22316 7100
rect 22340 7098 22396 7100
rect 22420 7098 22476 7100
rect 22500 7098 22556 7100
rect 22180 7046 22182 7098
rect 22182 7046 22234 7098
rect 22234 7046 22236 7098
rect 22260 7046 22298 7098
rect 22298 7046 22310 7098
rect 22310 7046 22316 7098
rect 22340 7046 22362 7098
rect 22362 7046 22374 7098
rect 22374 7046 22396 7098
rect 22420 7046 22426 7098
rect 22426 7046 22438 7098
rect 22438 7046 22476 7098
rect 22500 7046 22502 7098
rect 22502 7046 22554 7098
rect 22554 7046 22556 7098
rect 22180 7044 22236 7046
rect 22260 7044 22316 7046
rect 22340 7044 22396 7046
rect 22420 7044 22476 7046
rect 22500 7044 22556 7046
rect 28180 15802 28236 15804
rect 28260 15802 28316 15804
rect 28340 15802 28396 15804
rect 28420 15802 28476 15804
rect 28500 15802 28556 15804
rect 28180 15750 28182 15802
rect 28182 15750 28234 15802
rect 28234 15750 28236 15802
rect 28260 15750 28298 15802
rect 28298 15750 28310 15802
rect 28310 15750 28316 15802
rect 28340 15750 28362 15802
rect 28362 15750 28374 15802
rect 28374 15750 28396 15802
rect 28420 15750 28426 15802
rect 28426 15750 28438 15802
rect 28438 15750 28476 15802
rect 28500 15750 28502 15802
rect 28502 15750 28554 15802
rect 28554 15750 28556 15802
rect 28180 15748 28236 15750
rect 28260 15748 28316 15750
rect 28340 15748 28396 15750
rect 28420 15748 28476 15750
rect 28500 15748 28556 15750
rect 29090 16652 29146 16688
rect 29090 16632 29092 16652
rect 29092 16632 29144 16652
rect 29144 16632 29146 16652
rect 28920 16346 28976 16348
rect 29000 16346 29056 16348
rect 29080 16346 29136 16348
rect 29160 16346 29216 16348
rect 29240 16346 29296 16348
rect 28920 16294 28922 16346
rect 28922 16294 28974 16346
rect 28974 16294 28976 16346
rect 29000 16294 29038 16346
rect 29038 16294 29050 16346
rect 29050 16294 29056 16346
rect 29080 16294 29102 16346
rect 29102 16294 29114 16346
rect 29114 16294 29136 16346
rect 29160 16294 29166 16346
rect 29166 16294 29178 16346
rect 29178 16294 29216 16346
rect 29240 16294 29242 16346
rect 29242 16294 29294 16346
rect 29294 16294 29296 16346
rect 28920 16292 28976 16294
rect 29000 16292 29056 16294
rect 29080 16292 29136 16294
rect 29160 16292 29216 16294
rect 29240 16292 29296 16294
rect 28920 15258 28976 15260
rect 29000 15258 29056 15260
rect 29080 15258 29136 15260
rect 29160 15258 29216 15260
rect 29240 15258 29296 15260
rect 28920 15206 28922 15258
rect 28922 15206 28974 15258
rect 28974 15206 28976 15258
rect 29000 15206 29038 15258
rect 29038 15206 29050 15258
rect 29050 15206 29056 15258
rect 29080 15206 29102 15258
rect 29102 15206 29114 15258
rect 29114 15206 29136 15258
rect 29160 15206 29166 15258
rect 29166 15206 29178 15258
rect 29178 15206 29216 15258
rect 29240 15206 29242 15258
rect 29242 15206 29294 15258
rect 29294 15206 29296 15258
rect 28920 15204 28976 15206
rect 29000 15204 29056 15206
rect 29080 15204 29136 15206
rect 29160 15204 29216 15206
rect 29240 15204 29296 15206
rect 28180 14714 28236 14716
rect 28260 14714 28316 14716
rect 28340 14714 28396 14716
rect 28420 14714 28476 14716
rect 28500 14714 28556 14716
rect 28180 14662 28182 14714
rect 28182 14662 28234 14714
rect 28234 14662 28236 14714
rect 28260 14662 28298 14714
rect 28298 14662 28310 14714
rect 28310 14662 28316 14714
rect 28340 14662 28362 14714
rect 28362 14662 28374 14714
rect 28374 14662 28396 14714
rect 28420 14662 28426 14714
rect 28426 14662 28438 14714
rect 28438 14662 28476 14714
rect 28500 14662 28502 14714
rect 28502 14662 28554 14714
rect 28554 14662 28556 14714
rect 28180 14660 28236 14662
rect 28260 14660 28316 14662
rect 28340 14660 28396 14662
rect 28420 14660 28476 14662
rect 28500 14660 28556 14662
rect 28180 13626 28236 13628
rect 28260 13626 28316 13628
rect 28340 13626 28396 13628
rect 28420 13626 28476 13628
rect 28500 13626 28556 13628
rect 28180 13574 28182 13626
rect 28182 13574 28234 13626
rect 28234 13574 28236 13626
rect 28260 13574 28298 13626
rect 28298 13574 28310 13626
rect 28310 13574 28316 13626
rect 28340 13574 28362 13626
rect 28362 13574 28374 13626
rect 28374 13574 28396 13626
rect 28420 13574 28426 13626
rect 28426 13574 28438 13626
rect 28438 13574 28476 13626
rect 28500 13574 28502 13626
rect 28502 13574 28554 13626
rect 28554 13574 28556 13626
rect 28180 13572 28236 13574
rect 28260 13572 28316 13574
rect 28340 13572 28396 13574
rect 28420 13572 28476 13574
rect 28500 13572 28556 13574
rect 28920 14170 28976 14172
rect 29000 14170 29056 14172
rect 29080 14170 29136 14172
rect 29160 14170 29216 14172
rect 29240 14170 29296 14172
rect 28920 14118 28922 14170
rect 28922 14118 28974 14170
rect 28974 14118 28976 14170
rect 29000 14118 29038 14170
rect 29038 14118 29050 14170
rect 29050 14118 29056 14170
rect 29080 14118 29102 14170
rect 29102 14118 29114 14170
rect 29114 14118 29136 14170
rect 29160 14118 29166 14170
rect 29166 14118 29178 14170
rect 29178 14118 29216 14170
rect 29240 14118 29242 14170
rect 29242 14118 29294 14170
rect 29294 14118 29296 14170
rect 28920 14116 28976 14118
rect 29000 14116 29056 14118
rect 29080 14116 29136 14118
rect 29160 14116 29216 14118
rect 29240 14116 29296 14118
rect 28920 13082 28976 13084
rect 29000 13082 29056 13084
rect 29080 13082 29136 13084
rect 29160 13082 29216 13084
rect 29240 13082 29296 13084
rect 28920 13030 28922 13082
rect 28922 13030 28974 13082
rect 28974 13030 28976 13082
rect 29000 13030 29038 13082
rect 29038 13030 29050 13082
rect 29050 13030 29056 13082
rect 29080 13030 29102 13082
rect 29102 13030 29114 13082
rect 29114 13030 29136 13082
rect 29160 13030 29166 13082
rect 29166 13030 29178 13082
rect 29178 13030 29216 13082
rect 29240 13030 29242 13082
rect 29242 13030 29294 13082
rect 29294 13030 29296 13082
rect 28920 13028 28976 13030
rect 29000 13028 29056 13030
rect 29080 13028 29136 13030
rect 29160 13028 29216 13030
rect 29240 13028 29296 13030
rect 28180 12538 28236 12540
rect 28260 12538 28316 12540
rect 28340 12538 28396 12540
rect 28420 12538 28476 12540
rect 28500 12538 28556 12540
rect 28180 12486 28182 12538
rect 28182 12486 28234 12538
rect 28234 12486 28236 12538
rect 28260 12486 28298 12538
rect 28298 12486 28310 12538
rect 28310 12486 28316 12538
rect 28340 12486 28362 12538
rect 28362 12486 28374 12538
rect 28374 12486 28396 12538
rect 28420 12486 28426 12538
rect 28426 12486 28438 12538
rect 28438 12486 28476 12538
rect 28500 12486 28502 12538
rect 28502 12486 28554 12538
rect 28554 12486 28556 12538
rect 28180 12484 28236 12486
rect 28260 12484 28316 12486
rect 28340 12484 28396 12486
rect 28420 12484 28476 12486
rect 28500 12484 28556 12486
rect 22920 8730 22976 8732
rect 23000 8730 23056 8732
rect 23080 8730 23136 8732
rect 23160 8730 23216 8732
rect 23240 8730 23296 8732
rect 22920 8678 22922 8730
rect 22922 8678 22974 8730
rect 22974 8678 22976 8730
rect 23000 8678 23038 8730
rect 23038 8678 23050 8730
rect 23050 8678 23056 8730
rect 23080 8678 23102 8730
rect 23102 8678 23114 8730
rect 23114 8678 23136 8730
rect 23160 8678 23166 8730
rect 23166 8678 23178 8730
rect 23178 8678 23216 8730
rect 23240 8678 23242 8730
rect 23242 8678 23294 8730
rect 23294 8678 23296 8730
rect 22920 8676 22976 8678
rect 23000 8676 23056 8678
rect 23080 8676 23136 8678
rect 23160 8676 23216 8678
rect 23240 8676 23296 8678
rect 22920 7642 22976 7644
rect 23000 7642 23056 7644
rect 23080 7642 23136 7644
rect 23160 7642 23216 7644
rect 23240 7642 23296 7644
rect 22920 7590 22922 7642
rect 22922 7590 22974 7642
rect 22974 7590 22976 7642
rect 23000 7590 23038 7642
rect 23038 7590 23050 7642
rect 23050 7590 23056 7642
rect 23080 7590 23102 7642
rect 23102 7590 23114 7642
rect 23114 7590 23136 7642
rect 23160 7590 23166 7642
rect 23166 7590 23178 7642
rect 23178 7590 23216 7642
rect 23240 7590 23242 7642
rect 23242 7590 23294 7642
rect 23294 7590 23296 7642
rect 22920 7588 22976 7590
rect 23000 7588 23056 7590
rect 23080 7588 23136 7590
rect 23160 7588 23216 7590
rect 23240 7588 23296 7590
rect 22920 6554 22976 6556
rect 23000 6554 23056 6556
rect 23080 6554 23136 6556
rect 23160 6554 23216 6556
rect 23240 6554 23296 6556
rect 22920 6502 22922 6554
rect 22922 6502 22974 6554
rect 22974 6502 22976 6554
rect 23000 6502 23038 6554
rect 23038 6502 23050 6554
rect 23050 6502 23056 6554
rect 23080 6502 23102 6554
rect 23102 6502 23114 6554
rect 23114 6502 23136 6554
rect 23160 6502 23166 6554
rect 23166 6502 23178 6554
rect 23178 6502 23216 6554
rect 23240 6502 23242 6554
rect 23242 6502 23294 6554
rect 23294 6502 23296 6554
rect 22920 6500 22976 6502
rect 23000 6500 23056 6502
rect 23080 6500 23136 6502
rect 23160 6500 23216 6502
rect 23240 6500 23296 6502
rect 28920 11994 28976 11996
rect 29000 11994 29056 11996
rect 29080 11994 29136 11996
rect 29160 11994 29216 11996
rect 29240 11994 29296 11996
rect 28920 11942 28922 11994
rect 28922 11942 28974 11994
rect 28974 11942 28976 11994
rect 29000 11942 29038 11994
rect 29038 11942 29050 11994
rect 29050 11942 29056 11994
rect 29080 11942 29102 11994
rect 29102 11942 29114 11994
rect 29114 11942 29136 11994
rect 29160 11942 29166 11994
rect 29166 11942 29178 11994
rect 29178 11942 29216 11994
rect 29240 11942 29242 11994
rect 29242 11942 29294 11994
rect 29294 11942 29296 11994
rect 28920 11940 28976 11942
rect 29000 11940 29056 11942
rect 29080 11940 29136 11942
rect 29160 11940 29216 11942
rect 29240 11940 29296 11942
rect 28180 11450 28236 11452
rect 28260 11450 28316 11452
rect 28340 11450 28396 11452
rect 28420 11450 28476 11452
rect 28500 11450 28556 11452
rect 28180 11398 28182 11450
rect 28182 11398 28234 11450
rect 28234 11398 28236 11450
rect 28260 11398 28298 11450
rect 28298 11398 28310 11450
rect 28310 11398 28316 11450
rect 28340 11398 28362 11450
rect 28362 11398 28374 11450
rect 28374 11398 28396 11450
rect 28420 11398 28426 11450
rect 28426 11398 28438 11450
rect 28438 11398 28476 11450
rect 28500 11398 28502 11450
rect 28502 11398 28554 11450
rect 28554 11398 28556 11450
rect 28180 11396 28236 11398
rect 28260 11396 28316 11398
rect 28340 11396 28396 11398
rect 28420 11396 28476 11398
rect 28500 11396 28556 11398
rect 28920 10906 28976 10908
rect 29000 10906 29056 10908
rect 29080 10906 29136 10908
rect 29160 10906 29216 10908
rect 29240 10906 29296 10908
rect 28920 10854 28922 10906
rect 28922 10854 28974 10906
rect 28974 10854 28976 10906
rect 29000 10854 29038 10906
rect 29038 10854 29050 10906
rect 29050 10854 29056 10906
rect 29080 10854 29102 10906
rect 29102 10854 29114 10906
rect 29114 10854 29136 10906
rect 29160 10854 29166 10906
rect 29166 10854 29178 10906
rect 29178 10854 29216 10906
rect 29240 10854 29242 10906
rect 29242 10854 29294 10906
rect 29294 10854 29296 10906
rect 28920 10852 28976 10854
rect 29000 10852 29056 10854
rect 29080 10852 29136 10854
rect 29160 10852 29216 10854
rect 29240 10852 29296 10854
rect 22180 6010 22236 6012
rect 22260 6010 22316 6012
rect 22340 6010 22396 6012
rect 22420 6010 22476 6012
rect 22500 6010 22556 6012
rect 22180 5958 22182 6010
rect 22182 5958 22234 6010
rect 22234 5958 22236 6010
rect 22260 5958 22298 6010
rect 22298 5958 22310 6010
rect 22310 5958 22316 6010
rect 22340 5958 22362 6010
rect 22362 5958 22374 6010
rect 22374 5958 22396 6010
rect 22420 5958 22426 6010
rect 22426 5958 22438 6010
rect 22438 5958 22476 6010
rect 22500 5958 22502 6010
rect 22502 5958 22554 6010
rect 22554 5958 22556 6010
rect 22180 5956 22236 5958
rect 22260 5956 22316 5958
rect 22340 5956 22396 5958
rect 22420 5956 22476 5958
rect 22500 5956 22556 5958
rect 26882 8472 26938 8528
rect 28180 10362 28236 10364
rect 28260 10362 28316 10364
rect 28340 10362 28396 10364
rect 28420 10362 28476 10364
rect 28500 10362 28556 10364
rect 28180 10310 28182 10362
rect 28182 10310 28234 10362
rect 28234 10310 28236 10362
rect 28260 10310 28298 10362
rect 28298 10310 28310 10362
rect 28310 10310 28316 10362
rect 28340 10310 28362 10362
rect 28362 10310 28374 10362
rect 28374 10310 28396 10362
rect 28420 10310 28426 10362
rect 28426 10310 28438 10362
rect 28438 10310 28476 10362
rect 28500 10310 28502 10362
rect 28502 10310 28554 10362
rect 28554 10310 28556 10362
rect 28180 10308 28236 10310
rect 28260 10308 28316 10310
rect 28340 10308 28396 10310
rect 28420 10308 28476 10310
rect 28500 10308 28556 10310
rect 28920 9818 28976 9820
rect 29000 9818 29056 9820
rect 29080 9818 29136 9820
rect 29160 9818 29216 9820
rect 29240 9818 29296 9820
rect 28920 9766 28922 9818
rect 28922 9766 28974 9818
rect 28974 9766 28976 9818
rect 29000 9766 29038 9818
rect 29038 9766 29050 9818
rect 29050 9766 29056 9818
rect 29080 9766 29102 9818
rect 29102 9766 29114 9818
rect 29114 9766 29136 9818
rect 29160 9766 29166 9818
rect 29166 9766 29178 9818
rect 29178 9766 29216 9818
rect 29240 9766 29242 9818
rect 29242 9766 29294 9818
rect 29294 9766 29296 9818
rect 28920 9764 28976 9766
rect 29000 9764 29056 9766
rect 29080 9764 29136 9766
rect 29160 9764 29216 9766
rect 29240 9764 29296 9766
rect 28180 9274 28236 9276
rect 28260 9274 28316 9276
rect 28340 9274 28396 9276
rect 28420 9274 28476 9276
rect 28500 9274 28556 9276
rect 28180 9222 28182 9274
rect 28182 9222 28234 9274
rect 28234 9222 28236 9274
rect 28260 9222 28298 9274
rect 28298 9222 28310 9274
rect 28310 9222 28316 9274
rect 28340 9222 28362 9274
rect 28362 9222 28374 9274
rect 28374 9222 28396 9274
rect 28420 9222 28426 9274
rect 28426 9222 28438 9274
rect 28438 9222 28476 9274
rect 28500 9222 28502 9274
rect 28502 9222 28554 9274
rect 28554 9222 28556 9274
rect 28180 9220 28236 9222
rect 28260 9220 28316 9222
rect 28340 9220 28396 9222
rect 28420 9220 28476 9222
rect 28500 9220 28556 9222
rect 28180 8186 28236 8188
rect 28260 8186 28316 8188
rect 28340 8186 28396 8188
rect 28420 8186 28476 8188
rect 28500 8186 28556 8188
rect 28180 8134 28182 8186
rect 28182 8134 28234 8186
rect 28234 8134 28236 8186
rect 28260 8134 28298 8186
rect 28298 8134 28310 8186
rect 28310 8134 28316 8186
rect 28340 8134 28362 8186
rect 28362 8134 28374 8186
rect 28374 8134 28396 8186
rect 28420 8134 28426 8186
rect 28426 8134 28438 8186
rect 28438 8134 28476 8186
rect 28500 8134 28502 8186
rect 28502 8134 28554 8186
rect 28554 8134 28556 8186
rect 28180 8132 28236 8134
rect 28260 8132 28316 8134
rect 28340 8132 28396 8134
rect 28420 8132 28476 8134
rect 28500 8132 28556 8134
rect 30930 16632 30986 16688
rect 28920 8730 28976 8732
rect 29000 8730 29056 8732
rect 29080 8730 29136 8732
rect 29160 8730 29216 8732
rect 29240 8730 29296 8732
rect 28920 8678 28922 8730
rect 28922 8678 28974 8730
rect 28974 8678 28976 8730
rect 29000 8678 29038 8730
rect 29038 8678 29050 8730
rect 29050 8678 29056 8730
rect 29080 8678 29102 8730
rect 29102 8678 29114 8730
rect 29114 8678 29136 8730
rect 29160 8678 29166 8730
rect 29166 8678 29178 8730
rect 29178 8678 29216 8730
rect 29240 8678 29242 8730
rect 29242 8678 29294 8730
rect 29294 8678 29296 8730
rect 28920 8676 28976 8678
rect 29000 8676 29056 8678
rect 29080 8676 29136 8678
rect 29160 8676 29216 8678
rect 29240 8676 29296 8678
rect 28920 7642 28976 7644
rect 29000 7642 29056 7644
rect 29080 7642 29136 7644
rect 29160 7642 29216 7644
rect 29240 7642 29296 7644
rect 28920 7590 28922 7642
rect 28922 7590 28974 7642
rect 28974 7590 28976 7642
rect 29000 7590 29038 7642
rect 29038 7590 29050 7642
rect 29050 7590 29056 7642
rect 29080 7590 29102 7642
rect 29102 7590 29114 7642
rect 29114 7590 29136 7642
rect 29160 7590 29166 7642
rect 29166 7590 29178 7642
rect 29178 7590 29216 7642
rect 29240 7590 29242 7642
rect 29242 7590 29294 7642
rect 29294 7590 29296 7642
rect 28920 7588 28976 7590
rect 29000 7588 29056 7590
rect 29080 7588 29136 7590
rect 29160 7588 29216 7590
rect 29240 7588 29296 7590
rect 28180 7098 28236 7100
rect 28260 7098 28316 7100
rect 28340 7098 28396 7100
rect 28420 7098 28476 7100
rect 28500 7098 28556 7100
rect 28180 7046 28182 7098
rect 28182 7046 28234 7098
rect 28234 7046 28236 7098
rect 28260 7046 28298 7098
rect 28298 7046 28310 7098
rect 28310 7046 28316 7098
rect 28340 7046 28362 7098
rect 28362 7046 28374 7098
rect 28374 7046 28396 7098
rect 28420 7046 28426 7098
rect 28426 7046 28438 7098
rect 28438 7046 28476 7098
rect 28500 7046 28502 7098
rect 28502 7046 28554 7098
rect 28554 7046 28556 7098
rect 28180 7044 28236 7046
rect 28260 7044 28316 7046
rect 28340 7044 28396 7046
rect 28420 7044 28476 7046
rect 28500 7044 28556 7046
rect 28920 6554 28976 6556
rect 29000 6554 29056 6556
rect 29080 6554 29136 6556
rect 29160 6554 29216 6556
rect 29240 6554 29296 6556
rect 28920 6502 28922 6554
rect 28922 6502 28974 6554
rect 28974 6502 28976 6554
rect 29000 6502 29038 6554
rect 29038 6502 29050 6554
rect 29050 6502 29056 6554
rect 29080 6502 29102 6554
rect 29102 6502 29114 6554
rect 29114 6502 29136 6554
rect 29160 6502 29166 6554
rect 29166 6502 29178 6554
rect 29178 6502 29216 6554
rect 29240 6502 29242 6554
rect 29242 6502 29294 6554
rect 29294 6502 29296 6554
rect 28920 6500 28976 6502
rect 29000 6500 29056 6502
rect 29080 6500 29136 6502
rect 29160 6500 29216 6502
rect 29240 6500 29296 6502
rect 28180 6010 28236 6012
rect 28260 6010 28316 6012
rect 28340 6010 28396 6012
rect 28420 6010 28476 6012
rect 28500 6010 28556 6012
rect 28180 5958 28182 6010
rect 28182 5958 28234 6010
rect 28234 5958 28236 6010
rect 28260 5958 28298 6010
rect 28298 5958 28310 6010
rect 28310 5958 28316 6010
rect 28340 5958 28362 6010
rect 28362 5958 28374 6010
rect 28374 5958 28396 6010
rect 28420 5958 28426 6010
rect 28426 5958 28438 6010
rect 28438 5958 28476 6010
rect 28500 5958 28502 6010
rect 28502 5958 28554 6010
rect 28554 5958 28556 6010
rect 28180 5956 28236 5958
rect 28260 5956 28316 5958
rect 28340 5956 28396 5958
rect 28420 5956 28476 5958
rect 28500 5956 28556 5958
rect 22920 5466 22976 5468
rect 23000 5466 23056 5468
rect 23080 5466 23136 5468
rect 23160 5466 23216 5468
rect 23240 5466 23296 5468
rect 22920 5414 22922 5466
rect 22922 5414 22974 5466
rect 22974 5414 22976 5466
rect 23000 5414 23038 5466
rect 23038 5414 23050 5466
rect 23050 5414 23056 5466
rect 23080 5414 23102 5466
rect 23102 5414 23114 5466
rect 23114 5414 23136 5466
rect 23160 5414 23166 5466
rect 23166 5414 23178 5466
rect 23178 5414 23216 5466
rect 23240 5414 23242 5466
rect 23242 5414 23294 5466
rect 23294 5414 23296 5466
rect 22920 5412 22976 5414
rect 23000 5412 23056 5414
rect 23080 5412 23136 5414
rect 23160 5412 23216 5414
rect 23240 5412 23296 5414
rect 28920 5466 28976 5468
rect 29000 5466 29056 5468
rect 29080 5466 29136 5468
rect 29160 5466 29216 5468
rect 29240 5466 29296 5468
rect 28920 5414 28922 5466
rect 28922 5414 28974 5466
rect 28974 5414 28976 5466
rect 29000 5414 29038 5466
rect 29038 5414 29050 5466
rect 29050 5414 29056 5466
rect 29080 5414 29102 5466
rect 29102 5414 29114 5466
rect 29114 5414 29136 5466
rect 29160 5414 29166 5466
rect 29166 5414 29178 5466
rect 29178 5414 29216 5466
rect 29240 5414 29242 5466
rect 29242 5414 29294 5466
rect 29294 5414 29296 5466
rect 28920 5412 28976 5414
rect 29000 5412 29056 5414
rect 29080 5412 29136 5414
rect 29160 5412 29216 5414
rect 29240 5412 29296 5414
rect 22180 4922 22236 4924
rect 22260 4922 22316 4924
rect 22340 4922 22396 4924
rect 22420 4922 22476 4924
rect 22500 4922 22556 4924
rect 22180 4870 22182 4922
rect 22182 4870 22234 4922
rect 22234 4870 22236 4922
rect 22260 4870 22298 4922
rect 22298 4870 22310 4922
rect 22310 4870 22316 4922
rect 22340 4870 22362 4922
rect 22362 4870 22374 4922
rect 22374 4870 22396 4922
rect 22420 4870 22426 4922
rect 22426 4870 22438 4922
rect 22438 4870 22476 4922
rect 22500 4870 22502 4922
rect 22502 4870 22554 4922
rect 22554 4870 22556 4922
rect 22180 4868 22236 4870
rect 22260 4868 22316 4870
rect 22340 4868 22396 4870
rect 22420 4868 22476 4870
rect 22500 4868 22556 4870
rect 28180 4922 28236 4924
rect 28260 4922 28316 4924
rect 28340 4922 28396 4924
rect 28420 4922 28476 4924
rect 28500 4922 28556 4924
rect 28180 4870 28182 4922
rect 28182 4870 28234 4922
rect 28234 4870 28236 4922
rect 28260 4870 28298 4922
rect 28298 4870 28310 4922
rect 28310 4870 28316 4922
rect 28340 4870 28362 4922
rect 28362 4870 28374 4922
rect 28374 4870 28396 4922
rect 28420 4870 28426 4922
rect 28426 4870 28438 4922
rect 28438 4870 28476 4922
rect 28500 4870 28502 4922
rect 28502 4870 28554 4922
rect 28554 4870 28556 4922
rect 28180 4868 28236 4870
rect 28260 4868 28316 4870
rect 28340 4868 28396 4870
rect 28420 4868 28476 4870
rect 28500 4868 28556 4870
rect 16180 3834 16236 3836
rect 16260 3834 16316 3836
rect 16340 3834 16396 3836
rect 16420 3834 16476 3836
rect 16500 3834 16556 3836
rect 16180 3782 16182 3834
rect 16182 3782 16234 3834
rect 16234 3782 16236 3834
rect 16260 3782 16298 3834
rect 16298 3782 16310 3834
rect 16310 3782 16316 3834
rect 16340 3782 16362 3834
rect 16362 3782 16374 3834
rect 16374 3782 16396 3834
rect 16420 3782 16426 3834
rect 16426 3782 16438 3834
rect 16438 3782 16476 3834
rect 16500 3782 16502 3834
rect 16502 3782 16554 3834
rect 16554 3782 16556 3834
rect 16180 3780 16236 3782
rect 16260 3780 16316 3782
rect 16340 3780 16396 3782
rect 16420 3780 16476 3782
rect 16500 3780 16556 3782
rect 4180 2746 4236 2748
rect 4260 2746 4316 2748
rect 4340 2746 4396 2748
rect 4420 2746 4476 2748
rect 4500 2746 4556 2748
rect 4180 2694 4182 2746
rect 4182 2694 4234 2746
rect 4234 2694 4236 2746
rect 4260 2694 4298 2746
rect 4298 2694 4310 2746
rect 4310 2694 4316 2746
rect 4340 2694 4362 2746
rect 4362 2694 4374 2746
rect 4374 2694 4396 2746
rect 4420 2694 4426 2746
rect 4426 2694 4438 2746
rect 4438 2694 4476 2746
rect 4500 2694 4502 2746
rect 4502 2694 4554 2746
rect 4554 2694 4556 2746
rect 4180 2692 4236 2694
rect 4260 2692 4316 2694
rect 4340 2692 4396 2694
rect 4420 2692 4476 2694
rect 4500 2692 4556 2694
rect 10180 2746 10236 2748
rect 10260 2746 10316 2748
rect 10340 2746 10396 2748
rect 10420 2746 10476 2748
rect 10500 2746 10556 2748
rect 10180 2694 10182 2746
rect 10182 2694 10234 2746
rect 10234 2694 10236 2746
rect 10260 2694 10298 2746
rect 10298 2694 10310 2746
rect 10310 2694 10316 2746
rect 10340 2694 10362 2746
rect 10362 2694 10374 2746
rect 10374 2694 10396 2746
rect 10420 2694 10426 2746
rect 10426 2694 10438 2746
rect 10438 2694 10476 2746
rect 10500 2694 10502 2746
rect 10502 2694 10554 2746
rect 10554 2694 10556 2746
rect 10180 2692 10236 2694
rect 10260 2692 10316 2694
rect 10340 2692 10396 2694
rect 10420 2692 10476 2694
rect 10500 2692 10556 2694
rect 16920 4378 16976 4380
rect 17000 4378 17056 4380
rect 17080 4378 17136 4380
rect 17160 4378 17216 4380
rect 17240 4378 17296 4380
rect 16920 4326 16922 4378
rect 16922 4326 16974 4378
rect 16974 4326 16976 4378
rect 17000 4326 17038 4378
rect 17038 4326 17050 4378
rect 17050 4326 17056 4378
rect 17080 4326 17102 4378
rect 17102 4326 17114 4378
rect 17114 4326 17136 4378
rect 17160 4326 17166 4378
rect 17166 4326 17178 4378
rect 17178 4326 17216 4378
rect 17240 4326 17242 4378
rect 17242 4326 17294 4378
rect 17294 4326 17296 4378
rect 16920 4324 16976 4326
rect 17000 4324 17056 4326
rect 17080 4324 17136 4326
rect 17160 4324 17216 4326
rect 17240 4324 17296 4326
rect 22920 4378 22976 4380
rect 23000 4378 23056 4380
rect 23080 4378 23136 4380
rect 23160 4378 23216 4380
rect 23240 4378 23296 4380
rect 22920 4326 22922 4378
rect 22922 4326 22974 4378
rect 22974 4326 22976 4378
rect 23000 4326 23038 4378
rect 23038 4326 23050 4378
rect 23050 4326 23056 4378
rect 23080 4326 23102 4378
rect 23102 4326 23114 4378
rect 23114 4326 23136 4378
rect 23160 4326 23166 4378
rect 23166 4326 23178 4378
rect 23178 4326 23216 4378
rect 23240 4326 23242 4378
rect 23242 4326 23294 4378
rect 23294 4326 23296 4378
rect 22920 4324 22976 4326
rect 23000 4324 23056 4326
rect 23080 4324 23136 4326
rect 23160 4324 23216 4326
rect 23240 4324 23296 4326
rect 28920 4378 28976 4380
rect 29000 4378 29056 4380
rect 29080 4378 29136 4380
rect 29160 4378 29216 4380
rect 29240 4378 29296 4380
rect 28920 4326 28922 4378
rect 28922 4326 28974 4378
rect 28974 4326 28976 4378
rect 29000 4326 29038 4378
rect 29038 4326 29050 4378
rect 29050 4326 29056 4378
rect 29080 4326 29102 4378
rect 29102 4326 29114 4378
rect 29114 4326 29136 4378
rect 29160 4326 29166 4378
rect 29166 4326 29178 4378
rect 29178 4326 29216 4378
rect 29240 4326 29242 4378
rect 29242 4326 29294 4378
rect 29294 4326 29296 4378
rect 28920 4324 28976 4326
rect 29000 4324 29056 4326
rect 29080 4324 29136 4326
rect 29160 4324 29216 4326
rect 29240 4324 29296 4326
rect 22180 3834 22236 3836
rect 22260 3834 22316 3836
rect 22340 3834 22396 3836
rect 22420 3834 22476 3836
rect 22500 3834 22556 3836
rect 22180 3782 22182 3834
rect 22182 3782 22234 3834
rect 22234 3782 22236 3834
rect 22260 3782 22298 3834
rect 22298 3782 22310 3834
rect 22310 3782 22316 3834
rect 22340 3782 22362 3834
rect 22362 3782 22374 3834
rect 22374 3782 22396 3834
rect 22420 3782 22426 3834
rect 22426 3782 22438 3834
rect 22438 3782 22476 3834
rect 22500 3782 22502 3834
rect 22502 3782 22554 3834
rect 22554 3782 22556 3834
rect 22180 3780 22236 3782
rect 22260 3780 22316 3782
rect 22340 3780 22396 3782
rect 22420 3780 22476 3782
rect 22500 3780 22556 3782
rect 28180 3834 28236 3836
rect 28260 3834 28316 3836
rect 28340 3834 28396 3836
rect 28420 3834 28476 3836
rect 28500 3834 28556 3836
rect 28180 3782 28182 3834
rect 28182 3782 28234 3834
rect 28234 3782 28236 3834
rect 28260 3782 28298 3834
rect 28298 3782 28310 3834
rect 28310 3782 28316 3834
rect 28340 3782 28362 3834
rect 28362 3782 28374 3834
rect 28374 3782 28396 3834
rect 28420 3782 28426 3834
rect 28426 3782 28438 3834
rect 28438 3782 28476 3834
rect 28500 3782 28502 3834
rect 28502 3782 28554 3834
rect 28554 3782 28556 3834
rect 28180 3780 28236 3782
rect 28260 3780 28316 3782
rect 28340 3780 28396 3782
rect 28420 3780 28476 3782
rect 28500 3780 28556 3782
rect 16920 3290 16976 3292
rect 17000 3290 17056 3292
rect 17080 3290 17136 3292
rect 17160 3290 17216 3292
rect 17240 3290 17296 3292
rect 16920 3238 16922 3290
rect 16922 3238 16974 3290
rect 16974 3238 16976 3290
rect 17000 3238 17038 3290
rect 17038 3238 17050 3290
rect 17050 3238 17056 3290
rect 17080 3238 17102 3290
rect 17102 3238 17114 3290
rect 17114 3238 17136 3290
rect 17160 3238 17166 3290
rect 17166 3238 17178 3290
rect 17178 3238 17216 3290
rect 17240 3238 17242 3290
rect 17242 3238 17294 3290
rect 17294 3238 17296 3290
rect 16920 3236 16976 3238
rect 17000 3236 17056 3238
rect 17080 3236 17136 3238
rect 17160 3236 17216 3238
rect 17240 3236 17296 3238
rect 16180 2746 16236 2748
rect 16260 2746 16316 2748
rect 16340 2746 16396 2748
rect 16420 2746 16476 2748
rect 16500 2746 16556 2748
rect 16180 2694 16182 2746
rect 16182 2694 16234 2746
rect 16234 2694 16236 2746
rect 16260 2694 16298 2746
rect 16298 2694 16310 2746
rect 16310 2694 16316 2746
rect 16340 2694 16362 2746
rect 16362 2694 16374 2746
rect 16374 2694 16396 2746
rect 16420 2694 16426 2746
rect 16426 2694 16438 2746
rect 16438 2694 16476 2746
rect 16500 2694 16502 2746
rect 16502 2694 16554 2746
rect 16554 2694 16556 2746
rect 16180 2692 16236 2694
rect 16260 2692 16316 2694
rect 16340 2692 16396 2694
rect 16420 2692 16476 2694
rect 16500 2692 16556 2694
rect 17038 2488 17094 2544
rect 22920 3290 22976 3292
rect 23000 3290 23056 3292
rect 23080 3290 23136 3292
rect 23160 3290 23216 3292
rect 23240 3290 23296 3292
rect 22920 3238 22922 3290
rect 22922 3238 22974 3290
rect 22974 3238 22976 3290
rect 23000 3238 23038 3290
rect 23038 3238 23050 3290
rect 23050 3238 23056 3290
rect 23080 3238 23102 3290
rect 23102 3238 23114 3290
rect 23114 3238 23136 3290
rect 23160 3238 23166 3290
rect 23166 3238 23178 3290
rect 23178 3238 23216 3290
rect 23240 3238 23242 3290
rect 23242 3238 23294 3290
rect 23294 3238 23296 3290
rect 22920 3236 22976 3238
rect 23000 3236 23056 3238
rect 23080 3236 23136 3238
rect 23160 3236 23216 3238
rect 23240 3236 23296 3238
rect 28920 3290 28976 3292
rect 29000 3290 29056 3292
rect 29080 3290 29136 3292
rect 29160 3290 29216 3292
rect 29240 3290 29296 3292
rect 28920 3238 28922 3290
rect 28922 3238 28974 3290
rect 28974 3238 28976 3290
rect 29000 3238 29038 3290
rect 29038 3238 29050 3290
rect 29050 3238 29056 3290
rect 29080 3238 29102 3290
rect 29102 3238 29114 3290
rect 29114 3238 29136 3290
rect 29160 3238 29166 3290
rect 29166 3238 29178 3290
rect 29178 3238 29216 3290
rect 29240 3238 29242 3290
rect 29242 3238 29294 3290
rect 29294 3238 29296 3290
rect 28920 3236 28976 3238
rect 29000 3236 29056 3238
rect 29080 3236 29136 3238
rect 29160 3236 29216 3238
rect 29240 3236 29296 3238
rect 22180 2746 22236 2748
rect 22260 2746 22316 2748
rect 22340 2746 22396 2748
rect 22420 2746 22476 2748
rect 22500 2746 22556 2748
rect 22180 2694 22182 2746
rect 22182 2694 22234 2746
rect 22234 2694 22236 2746
rect 22260 2694 22298 2746
rect 22298 2694 22310 2746
rect 22310 2694 22316 2746
rect 22340 2694 22362 2746
rect 22362 2694 22374 2746
rect 22374 2694 22396 2746
rect 22420 2694 22426 2746
rect 22426 2694 22438 2746
rect 22438 2694 22476 2746
rect 22500 2694 22502 2746
rect 22502 2694 22554 2746
rect 22554 2694 22556 2746
rect 22180 2692 22236 2694
rect 22260 2692 22316 2694
rect 22340 2692 22396 2694
rect 22420 2692 22476 2694
rect 22500 2692 22556 2694
rect 28180 2746 28236 2748
rect 28260 2746 28316 2748
rect 28340 2746 28396 2748
rect 28420 2746 28476 2748
rect 28500 2746 28556 2748
rect 28180 2694 28182 2746
rect 28182 2694 28234 2746
rect 28234 2694 28236 2746
rect 28260 2694 28298 2746
rect 28298 2694 28310 2746
rect 28310 2694 28316 2746
rect 28340 2694 28362 2746
rect 28362 2694 28374 2746
rect 28374 2694 28396 2746
rect 28420 2694 28426 2746
rect 28426 2694 28438 2746
rect 28438 2694 28476 2746
rect 28500 2694 28502 2746
rect 28502 2694 28554 2746
rect 28554 2694 28556 2746
rect 28180 2692 28236 2694
rect 28260 2692 28316 2694
rect 28340 2692 28396 2694
rect 28420 2692 28476 2694
rect 28500 2692 28556 2694
rect 31850 19760 31906 19816
rect 31482 13640 31538 13696
rect 31850 7520 31906 7576
rect 4920 2202 4976 2204
rect 5000 2202 5056 2204
rect 5080 2202 5136 2204
rect 5160 2202 5216 2204
rect 5240 2202 5296 2204
rect 4920 2150 4922 2202
rect 4922 2150 4974 2202
rect 4974 2150 4976 2202
rect 5000 2150 5038 2202
rect 5038 2150 5050 2202
rect 5050 2150 5056 2202
rect 5080 2150 5102 2202
rect 5102 2150 5114 2202
rect 5114 2150 5136 2202
rect 5160 2150 5166 2202
rect 5166 2150 5178 2202
rect 5178 2150 5216 2202
rect 5240 2150 5242 2202
rect 5242 2150 5294 2202
rect 5294 2150 5296 2202
rect 4920 2148 4976 2150
rect 5000 2148 5056 2150
rect 5080 2148 5136 2150
rect 5160 2148 5216 2150
rect 5240 2148 5296 2150
rect 10920 2202 10976 2204
rect 11000 2202 11056 2204
rect 11080 2202 11136 2204
rect 11160 2202 11216 2204
rect 11240 2202 11296 2204
rect 10920 2150 10922 2202
rect 10922 2150 10974 2202
rect 10974 2150 10976 2202
rect 11000 2150 11038 2202
rect 11038 2150 11050 2202
rect 11050 2150 11056 2202
rect 11080 2150 11102 2202
rect 11102 2150 11114 2202
rect 11114 2150 11136 2202
rect 11160 2150 11166 2202
rect 11166 2150 11178 2202
rect 11178 2150 11216 2202
rect 11240 2150 11242 2202
rect 11242 2150 11294 2202
rect 11294 2150 11296 2202
rect 10920 2148 10976 2150
rect 11000 2148 11056 2150
rect 11080 2148 11136 2150
rect 11160 2148 11216 2150
rect 11240 2148 11296 2150
rect 16920 2202 16976 2204
rect 17000 2202 17056 2204
rect 17080 2202 17136 2204
rect 17160 2202 17216 2204
rect 17240 2202 17296 2204
rect 16920 2150 16922 2202
rect 16922 2150 16974 2202
rect 16974 2150 16976 2202
rect 17000 2150 17038 2202
rect 17038 2150 17050 2202
rect 17050 2150 17056 2202
rect 17080 2150 17102 2202
rect 17102 2150 17114 2202
rect 17114 2150 17136 2202
rect 17160 2150 17166 2202
rect 17166 2150 17178 2202
rect 17178 2150 17216 2202
rect 17240 2150 17242 2202
rect 17242 2150 17294 2202
rect 17294 2150 17296 2202
rect 16920 2148 16976 2150
rect 17000 2148 17056 2150
rect 17080 2148 17136 2150
rect 17160 2148 17216 2150
rect 17240 2148 17296 2150
rect 22920 2202 22976 2204
rect 23000 2202 23056 2204
rect 23080 2202 23136 2204
rect 23160 2202 23216 2204
rect 23240 2202 23296 2204
rect 22920 2150 22922 2202
rect 22922 2150 22974 2202
rect 22974 2150 22976 2202
rect 23000 2150 23038 2202
rect 23038 2150 23050 2202
rect 23050 2150 23056 2202
rect 23080 2150 23102 2202
rect 23102 2150 23114 2202
rect 23114 2150 23136 2202
rect 23160 2150 23166 2202
rect 23166 2150 23178 2202
rect 23178 2150 23216 2202
rect 23240 2150 23242 2202
rect 23242 2150 23294 2202
rect 23294 2150 23296 2202
rect 22920 2148 22976 2150
rect 23000 2148 23056 2150
rect 23080 2148 23136 2150
rect 23160 2148 23216 2150
rect 23240 2148 23296 2150
rect 28920 2202 28976 2204
rect 29000 2202 29056 2204
rect 29080 2202 29136 2204
rect 29160 2202 29216 2204
rect 29240 2202 29296 2204
rect 28920 2150 28922 2202
rect 28922 2150 28974 2202
rect 28974 2150 28976 2202
rect 29000 2150 29038 2202
rect 29038 2150 29050 2202
rect 29050 2150 29056 2202
rect 29080 2150 29102 2202
rect 29102 2150 29114 2202
rect 29114 2150 29136 2202
rect 29160 2150 29166 2202
rect 29166 2150 29178 2202
rect 29178 2150 29216 2202
rect 29240 2150 29242 2202
rect 29242 2150 29294 2202
rect 29294 2150 29296 2202
rect 28920 2148 28976 2150
rect 29000 2148 29056 2150
rect 29080 2148 29136 2150
rect 29160 2148 29216 2150
rect 29240 2148 29296 2150
rect 31390 1400 31446 1456
<< metal3 >>
rect 4910 32672 5306 32673
rect 4910 32608 4916 32672
rect 4980 32608 4996 32672
rect 5060 32608 5076 32672
rect 5140 32608 5156 32672
rect 5220 32608 5236 32672
rect 5300 32608 5306 32672
rect 4910 32607 5306 32608
rect 10910 32672 11306 32673
rect 10910 32608 10916 32672
rect 10980 32608 10996 32672
rect 11060 32608 11076 32672
rect 11140 32608 11156 32672
rect 11220 32608 11236 32672
rect 11300 32608 11306 32672
rect 10910 32607 11306 32608
rect 16910 32672 17306 32673
rect 16910 32608 16916 32672
rect 16980 32608 16996 32672
rect 17060 32608 17076 32672
rect 17140 32608 17156 32672
rect 17220 32608 17236 32672
rect 17300 32608 17306 32672
rect 16910 32607 17306 32608
rect 22910 32672 23306 32673
rect 22910 32608 22916 32672
rect 22980 32608 22996 32672
rect 23060 32608 23076 32672
rect 23140 32608 23156 32672
rect 23220 32608 23236 32672
rect 23300 32608 23306 32672
rect 22910 32607 23306 32608
rect 28910 32672 29306 32673
rect 28910 32608 28916 32672
rect 28980 32608 28996 32672
rect 29060 32608 29076 32672
rect 29140 32608 29156 32672
rect 29220 32608 29236 32672
rect 29300 32608 29306 32672
rect 28910 32607 29306 32608
rect 4170 32128 4566 32129
rect 4170 32064 4176 32128
rect 4240 32064 4256 32128
rect 4320 32064 4336 32128
rect 4400 32064 4416 32128
rect 4480 32064 4496 32128
rect 4560 32064 4566 32128
rect 4170 32063 4566 32064
rect 10170 32128 10566 32129
rect 10170 32064 10176 32128
rect 10240 32064 10256 32128
rect 10320 32064 10336 32128
rect 10400 32064 10416 32128
rect 10480 32064 10496 32128
rect 10560 32064 10566 32128
rect 10170 32063 10566 32064
rect 16170 32128 16566 32129
rect 16170 32064 16176 32128
rect 16240 32064 16256 32128
rect 16320 32064 16336 32128
rect 16400 32064 16416 32128
rect 16480 32064 16496 32128
rect 16560 32064 16566 32128
rect 16170 32063 16566 32064
rect 22170 32128 22566 32129
rect 22170 32064 22176 32128
rect 22240 32064 22256 32128
rect 22320 32064 22336 32128
rect 22400 32064 22416 32128
rect 22480 32064 22496 32128
rect 22560 32064 22566 32128
rect 22170 32063 22566 32064
rect 28170 32128 28566 32129
rect 28170 32064 28176 32128
rect 28240 32064 28256 32128
rect 28320 32064 28336 32128
rect 28400 32064 28416 32128
rect 28480 32064 28496 32128
rect 28560 32064 28566 32128
rect 28170 32063 28566 32064
rect 32174 32058 32974 32088
rect 28766 31998 32974 32058
rect 27838 31860 27844 31924
rect 27908 31922 27914 31924
rect 28766 31922 28826 31998
rect 32174 31968 32974 31998
rect 27908 31862 28826 31922
rect 27908 31860 27914 31862
rect 4910 31584 5306 31585
rect 4910 31520 4916 31584
rect 4980 31520 4996 31584
rect 5060 31520 5076 31584
rect 5140 31520 5156 31584
rect 5220 31520 5236 31584
rect 5300 31520 5306 31584
rect 4910 31519 5306 31520
rect 10910 31584 11306 31585
rect 10910 31520 10916 31584
rect 10980 31520 10996 31584
rect 11060 31520 11076 31584
rect 11140 31520 11156 31584
rect 11220 31520 11236 31584
rect 11300 31520 11306 31584
rect 10910 31519 11306 31520
rect 16910 31584 17306 31585
rect 16910 31520 16916 31584
rect 16980 31520 16996 31584
rect 17060 31520 17076 31584
rect 17140 31520 17156 31584
rect 17220 31520 17236 31584
rect 17300 31520 17306 31584
rect 16910 31519 17306 31520
rect 22910 31584 23306 31585
rect 22910 31520 22916 31584
rect 22980 31520 22996 31584
rect 23060 31520 23076 31584
rect 23140 31520 23156 31584
rect 23220 31520 23236 31584
rect 23300 31520 23306 31584
rect 22910 31519 23306 31520
rect 28910 31584 29306 31585
rect 28910 31520 28916 31584
rect 28980 31520 28996 31584
rect 29060 31520 29076 31584
rect 29140 31520 29156 31584
rect 29220 31520 29236 31584
rect 29300 31520 29306 31584
rect 28910 31519 29306 31520
rect 4170 31040 4566 31041
rect 4170 30976 4176 31040
rect 4240 30976 4256 31040
rect 4320 30976 4336 31040
rect 4400 30976 4416 31040
rect 4480 30976 4496 31040
rect 4560 30976 4566 31040
rect 4170 30975 4566 30976
rect 10170 31040 10566 31041
rect 10170 30976 10176 31040
rect 10240 30976 10256 31040
rect 10320 30976 10336 31040
rect 10400 30976 10416 31040
rect 10480 30976 10496 31040
rect 10560 30976 10566 31040
rect 10170 30975 10566 30976
rect 16170 31040 16566 31041
rect 16170 30976 16176 31040
rect 16240 30976 16256 31040
rect 16320 30976 16336 31040
rect 16400 30976 16416 31040
rect 16480 30976 16496 31040
rect 16560 30976 16566 31040
rect 16170 30975 16566 30976
rect 22170 31040 22566 31041
rect 22170 30976 22176 31040
rect 22240 30976 22256 31040
rect 22320 30976 22336 31040
rect 22400 30976 22416 31040
rect 22480 30976 22496 31040
rect 22560 30976 22566 31040
rect 22170 30975 22566 30976
rect 28170 31040 28566 31041
rect 28170 30976 28176 31040
rect 28240 30976 28256 31040
rect 28320 30976 28336 31040
rect 28400 30976 28416 31040
rect 28480 30976 28496 31040
rect 28560 30976 28566 31040
rect 28170 30975 28566 30976
rect 0 30698 800 30728
rect 933 30698 999 30701
rect 0 30696 999 30698
rect 0 30640 938 30696
rect 994 30640 999 30696
rect 0 30638 999 30640
rect 0 30608 800 30638
rect 933 30635 999 30638
rect 4910 30496 5306 30497
rect 4910 30432 4916 30496
rect 4980 30432 4996 30496
rect 5060 30432 5076 30496
rect 5140 30432 5156 30496
rect 5220 30432 5236 30496
rect 5300 30432 5306 30496
rect 4910 30431 5306 30432
rect 10910 30496 11306 30497
rect 10910 30432 10916 30496
rect 10980 30432 10996 30496
rect 11060 30432 11076 30496
rect 11140 30432 11156 30496
rect 11220 30432 11236 30496
rect 11300 30432 11306 30496
rect 10910 30431 11306 30432
rect 16910 30496 17306 30497
rect 16910 30432 16916 30496
rect 16980 30432 16996 30496
rect 17060 30432 17076 30496
rect 17140 30432 17156 30496
rect 17220 30432 17236 30496
rect 17300 30432 17306 30496
rect 16910 30431 17306 30432
rect 22910 30496 23306 30497
rect 22910 30432 22916 30496
rect 22980 30432 22996 30496
rect 23060 30432 23076 30496
rect 23140 30432 23156 30496
rect 23220 30432 23236 30496
rect 23300 30432 23306 30496
rect 22910 30431 23306 30432
rect 28910 30496 29306 30497
rect 28910 30432 28916 30496
rect 28980 30432 28996 30496
rect 29060 30432 29076 30496
rect 29140 30432 29156 30496
rect 29220 30432 29236 30496
rect 29300 30432 29306 30496
rect 28910 30431 29306 30432
rect 4170 29952 4566 29953
rect 4170 29888 4176 29952
rect 4240 29888 4256 29952
rect 4320 29888 4336 29952
rect 4400 29888 4416 29952
rect 4480 29888 4496 29952
rect 4560 29888 4566 29952
rect 4170 29887 4566 29888
rect 10170 29952 10566 29953
rect 10170 29888 10176 29952
rect 10240 29888 10256 29952
rect 10320 29888 10336 29952
rect 10400 29888 10416 29952
rect 10480 29888 10496 29952
rect 10560 29888 10566 29952
rect 10170 29887 10566 29888
rect 16170 29952 16566 29953
rect 16170 29888 16176 29952
rect 16240 29888 16256 29952
rect 16320 29888 16336 29952
rect 16400 29888 16416 29952
rect 16480 29888 16496 29952
rect 16560 29888 16566 29952
rect 16170 29887 16566 29888
rect 22170 29952 22566 29953
rect 22170 29888 22176 29952
rect 22240 29888 22256 29952
rect 22320 29888 22336 29952
rect 22400 29888 22416 29952
rect 22480 29888 22496 29952
rect 22560 29888 22566 29952
rect 22170 29887 22566 29888
rect 28170 29952 28566 29953
rect 28170 29888 28176 29952
rect 28240 29888 28256 29952
rect 28320 29888 28336 29952
rect 28400 29888 28416 29952
rect 28480 29888 28496 29952
rect 28560 29888 28566 29952
rect 28170 29887 28566 29888
rect 4910 29408 5306 29409
rect 4910 29344 4916 29408
rect 4980 29344 4996 29408
rect 5060 29344 5076 29408
rect 5140 29344 5156 29408
rect 5220 29344 5236 29408
rect 5300 29344 5306 29408
rect 4910 29343 5306 29344
rect 10910 29408 11306 29409
rect 10910 29344 10916 29408
rect 10980 29344 10996 29408
rect 11060 29344 11076 29408
rect 11140 29344 11156 29408
rect 11220 29344 11236 29408
rect 11300 29344 11306 29408
rect 10910 29343 11306 29344
rect 16910 29408 17306 29409
rect 16910 29344 16916 29408
rect 16980 29344 16996 29408
rect 17060 29344 17076 29408
rect 17140 29344 17156 29408
rect 17220 29344 17236 29408
rect 17300 29344 17306 29408
rect 16910 29343 17306 29344
rect 22910 29408 23306 29409
rect 22910 29344 22916 29408
rect 22980 29344 22996 29408
rect 23060 29344 23076 29408
rect 23140 29344 23156 29408
rect 23220 29344 23236 29408
rect 23300 29344 23306 29408
rect 22910 29343 23306 29344
rect 28910 29408 29306 29409
rect 28910 29344 28916 29408
rect 28980 29344 28996 29408
rect 29060 29344 29076 29408
rect 29140 29344 29156 29408
rect 29220 29344 29236 29408
rect 29300 29344 29306 29408
rect 28910 29343 29306 29344
rect 13997 29068 14063 29069
rect 13997 29066 14044 29068
rect 13952 29064 14044 29066
rect 13952 29008 14002 29064
rect 13952 29006 14044 29008
rect 13997 29004 14044 29006
rect 14108 29004 14114 29068
rect 13997 29003 14063 29004
rect 4170 28864 4566 28865
rect 4170 28800 4176 28864
rect 4240 28800 4256 28864
rect 4320 28800 4336 28864
rect 4400 28800 4416 28864
rect 4480 28800 4496 28864
rect 4560 28800 4566 28864
rect 4170 28799 4566 28800
rect 10170 28864 10566 28865
rect 10170 28800 10176 28864
rect 10240 28800 10256 28864
rect 10320 28800 10336 28864
rect 10400 28800 10416 28864
rect 10480 28800 10496 28864
rect 10560 28800 10566 28864
rect 10170 28799 10566 28800
rect 16170 28864 16566 28865
rect 16170 28800 16176 28864
rect 16240 28800 16256 28864
rect 16320 28800 16336 28864
rect 16400 28800 16416 28864
rect 16480 28800 16496 28864
rect 16560 28800 16566 28864
rect 16170 28799 16566 28800
rect 22170 28864 22566 28865
rect 22170 28800 22176 28864
rect 22240 28800 22256 28864
rect 22320 28800 22336 28864
rect 22400 28800 22416 28864
rect 22480 28800 22496 28864
rect 22560 28800 22566 28864
rect 22170 28799 22566 28800
rect 28170 28864 28566 28865
rect 28170 28800 28176 28864
rect 28240 28800 28256 28864
rect 28320 28800 28336 28864
rect 28400 28800 28416 28864
rect 28480 28800 28496 28864
rect 28560 28800 28566 28864
rect 28170 28799 28566 28800
rect 4910 28320 5306 28321
rect 4910 28256 4916 28320
rect 4980 28256 4996 28320
rect 5060 28256 5076 28320
rect 5140 28256 5156 28320
rect 5220 28256 5236 28320
rect 5300 28256 5306 28320
rect 4910 28255 5306 28256
rect 10910 28320 11306 28321
rect 10910 28256 10916 28320
rect 10980 28256 10996 28320
rect 11060 28256 11076 28320
rect 11140 28256 11156 28320
rect 11220 28256 11236 28320
rect 11300 28256 11306 28320
rect 10910 28255 11306 28256
rect 16910 28320 17306 28321
rect 16910 28256 16916 28320
rect 16980 28256 16996 28320
rect 17060 28256 17076 28320
rect 17140 28256 17156 28320
rect 17220 28256 17236 28320
rect 17300 28256 17306 28320
rect 16910 28255 17306 28256
rect 22910 28320 23306 28321
rect 22910 28256 22916 28320
rect 22980 28256 22996 28320
rect 23060 28256 23076 28320
rect 23140 28256 23156 28320
rect 23220 28256 23236 28320
rect 23300 28256 23306 28320
rect 22910 28255 23306 28256
rect 28910 28320 29306 28321
rect 28910 28256 28916 28320
rect 28980 28256 28996 28320
rect 29060 28256 29076 28320
rect 29140 28256 29156 28320
rect 29220 28256 29236 28320
rect 29300 28256 29306 28320
rect 28910 28255 29306 28256
rect 4170 27776 4566 27777
rect 4170 27712 4176 27776
rect 4240 27712 4256 27776
rect 4320 27712 4336 27776
rect 4400 27712 4416 27776
rect 4480 27712 4496 27776
rect 4560 27712 4566 27776
rect 4170 27711 4566 27712
rect 10170 27776 10566 27777
rect 10170 27712 10176 27776
rect 10240 27712 10256 27776
rect 10320 27712 10336 27776
rect 10400 27712 10416 27776
rect 10480 27712 10496 27776
rect 10560 27712 10566 27776
rect 10170 27711 10566 27712
rect 16170 27776 16566 27777
rect 16170 27712 16176 27776
rect 16240 27712 16256 27776
rect 16320 27712 16336 27776
rect 16400 27712 16416 27776
rect 16480 27712 16496 27776
rect 16560 27712 16566 27776
rect 16170 27711 16566 27712
rect 22170 27776 22566 27777
rect 22170 27712 22176 27776
rect 22240 27712 22256 27776
rect 22320 27712 22336 27776
rect 22400 27712 22416 27776
rect 22480 27712 22496 27776
rect 22560 27712 22566 27776
rect 22170 27711 22566 27712
rect 28170 27776 28566 27777
rect 28170 27712 28176 27776
rect 28240 27712 28256 27776
rect 28320 27712 28336 27776
rect 28400 27712 28416 27776
rect 28480 27712 28496 27776
rect 28560 27712 28566 27776
rect 28170 27711 28566 27712
rect 15929 27434 15995 27437
rect 17769 27434 17835 27437
rect 15929 27432 17835 27434
rect 15929 27376 15934 27432
rect 15990 27376 17774 27432
rect 17830 27376 17835 27432
rect 15929 27374 17835 27376
rect 15929 27371 15995 27374
rect 17769 27371 17835 27374
rect 4910 27232 5306 27233
rect 4910 27168 4916 27232
rect 4980 27168 4996 27232
rect 5060 27168 5076 27232
rect 5140 27168 5156 27232
rect 5220 27168 5236 27232
rect 5300 27168 5306 27232
rect 4910 27167 5306 27168
rect 10910 27232 11306 27233
rect 10910 27168 10916 27232
rect 10980 27168 10996 27232
rect 11060 27168 11076 27232
rect 11140 27168 11156 27232
rect 11220 27168 11236 27232
rect 11300 27168 11306 27232
rect 10910 27167 11306 27168
rect 16910 27232 17306 27233
rect 16910 27168 16916 27232
rect 16980 27168 16996 27232
rect 17060 27168 17076 27232
rect 17140 27168 17156 27232
rect 17220 27168 17236 27232
rect 17300 27168 17306 27232
rect 16910 27167 17306 27168
rect 22910 27232 23306 27233
rect 22910 27168 22916 27232
rect 22980 27168 22996 27232
rect 23060 27168 23076 27232
rect 23140 27168 23156 27232
rect 23220 27168 23236 27232
rect 23300 27168 23306 27232
rect 22910 27167 23306 27168
rect 28910 27232 29306 27233
rect 28910 27168 28916 27232
rect 28980 27168 28996 27232
rect 29060 27168 29076 27232
rect 29140 27168 29156 27232
rect 29220 27168 29236 27232
rect 29300 27168 29306 27232
rect 28910 27167 29306 27168
rect 9213 27026 9279 27029
rect 23749 27026 23815 27029
rect 9213 27024 23815 27026
rect 9213 26968 9218 27024
rect 9274 26968 23754 27024
rect 23810 26968 23815 27024
rect 9213 26966 23815 26968
rect 9213 26963 9279 26966
rect 23749 26963 23815 26966
rect 16113 26890 16179 26893
rect 17125 26890 17191 26893
rect 18045 26890 18111 26893
rect 16113 26888 18111 26890
rect 16113 26832 16118 26888
rect 16174 26832 17130 26888
rect 17186 26832 18050 26888
rect 18106 26832 18111 26888
rect 16113 26830 18111 26832
rect 16113 26827 16179 26830
rect 17125 26827 17191 26830
rect 18045 26827 18111 26830
rect 16849 26754 16915 26757
rect 18321 26754 18387 26757
rect 16849 26752 18387 26754
rect 16849 26696 16854 26752
rect 16910 26696 18326 26752
rect 18382 26696 18387 26752
rect 16849 26694 18387 26696
rect 16849 26691 16915 26694
rect 18321 26691 18387 26694
rect 4170 26688 4566 26689
rect 4170 26624 4176 26688
rect 4240 26624 4256 26688
rect 4320 26624 4336 26688
rect 4400 26624 4416 26688
rect 4480 26624 4496 26688
rect 4560 26624 4566 26688
rect 4170 26623 4566 26624
rect 10170 26688 10566 26689
rect 10170 26624 10176 26688
rect 10240 26624 10256 26688
rect 10320 26624 10336 26688
rect 10400 26624 10416 26688
rect 10480 26624 10496 26688
rect 10560 26624 10566 26688
rect 10170 26623 10566 26624
rect 16170 26688 16566 26689
rect 16170 26624 16176 26688
rect 16240 26624 16256 26688
rect 16320 26624 16336 26688
rect 16400 26624 16416 26688
rect 16480 26624 16496 26688
rect 16560 26624 16566 26688
rect 16170 26623 16566 26624
rect 22170 26688 22566 26689
rect 22170 26624 22176 26688
rect 22240 26624 22256 26688
rect 22320 26624 22336 26688
rect 22400 26624 22416 26688
rect 22480 26624 22496 26688
rect 22560 26624 22566 26688
rect 22170 26623 22566 26624
rect 28170 26688 28566 26689
rect 28170 26624 28176 26688
rect 28240 26624 28256 26688
rect 28320 26624 28336 26688
rect 28400 26624 28416 26688
rect 28480 26624 28496 26688
rect 28560 26624 28566 26688
rect 28170 26623 28566 26624
rect 4910 26144 5306 26145
rect 4910 26080 4916 26144
rect 4980 26080 4996 26144
rect 5060 26080 5076 26144
rect 5140 26080 5156 26144
rect 5220 26080 5236 26144
rect 5300 26080 5306 26144
rect 4910 26079 5306 26080
rect 10910 26144 11306 26145
rect 10910 26080 10916 26144
rect 10980 26080 10996 26144
rect 11060 26080 11076 26144
rect 11140 26080 11156 26144
rect 11220 26080 11236 26144
rect 11300 26080 11306 26144
rect 10910 26079 11306 26080
rect 16910 26144 17306 26145
rect 16910 26080 16916 26144
rect 16980 26080 16996 26144
rect 17060 26080 17076 26144
rect 17140 26080 17156 26144
rect 17220 26080 17236 26144
rect 17300 26080 17306 26144
rect 16910 26079 17306 26080
rect 22910 26144 23306 26145
rect 22910 26080 22916 26144
rect 22980 26080 22996 26144
rect 23060 26080 23076 26144
rect 23140 26080 23156 26144
rect 23220 26080 23236 26144
rect 23300 26080 23306 26144
rect 22910 26079 23306 26080
rect 28910 26144 29306 26145
rect 28910 26080 28916 26144
rect 28980 26080 28996 26144
rect 29060 26080 29076 26144
rect 29140 26080 29156 26144
rect 29220 26080 29236 26144
rect 29300 26080 29306 26144
rect 28910 26079 29306 26080
rect 31477 25938 31543 25941
rect 32174 25938 32974 25968
rect 31477 25936 32974 25938
rect 31477 25880 31482 25936
rect 31538 25880 32974 25936
rect 31477 25878 32974 25880
rect 31477 25875 31543 25878
rect 32174 25848 32974 25878
rect 4170 25600 4566 25601
rect 4170 25536 4176 25600
rect 4240 25536 4256 25600
rect 4320 25536 4336 25600
rect 4400 25536 4416 25600
rect 4480 25536 4496 25600
rect 4560 25536 4566 25600
rect 4170 25535 4566 25536
rect 10170 25600 10566 25601
rect 10170 25536 10176 25600
rect 10240 25536 10256 25600
rect 10320 25536 10336 25600
rect 10400 25536 10416 25600
rect 10480 25536 10496 25600
rect 10560 25536 10566 25600
rect 10170 25535 10566 25536
rect 16170 25600 16566 25601
rect 16170 25536 16176 25600
rect 16240 25536 16256 25600
rect 16320 25536 16336 25600
rect 16400 25536 16416 25600
rect 16480 25536 16496 25600
rect 16560 25536 16566 25600
rect 16170 25535 16566 25536
rect 22170 25600 22566 25601
rect 22170 25536 22176 25600
rect 22240 25536 22256 25600
rect 22320 25536 22336 25600
rect 22400 25536 22416 25600
rect 22480 25536 22496 25600
rect 22560 25536 22566 25600
rect 22170 25535 22566 25536
rect 28170 25600 28566 25601
rect 28170 25536 28176 25600
rect 28240 25536 28256 25600
rect 28320 25536 28336 25600
rect 28400 25536 28416 25600
rect 28480 25536 28496 25600
rect 28560 25536 28566 25600
rect 28170 25535 28566 25536
rect 4910 25056 5306 25057
rect 4910 24992 4916 25056
rect 4980 24992 4996 25056
rect 5060 24992 5076 25056
rect 5140 24992 5156 25056
rect 5220 24992 5236 25056
rect 5300 24992 5306 25056
rect 4910 24991 5306 24992
rect 10910 25056 11306 25057
rect 10910 24992 10916 25056
rect 10980 24992 10996 25056
rect 11060 24992 11076 25056
rect 11140 24992 11156 25056
rect 11220 24992 11236 25056
rect 11300 24992 11306 25056
rect 10910 24991 11306 24992
rect 16910 25056 17306 25057
rect 16910 24992 16916 25056
rect 16980 24992 16996 25056
rect 17060 24992 17076 25056
rect 17140 24992 17156 25056
rect 17220 24992 17236 25056
rect 17300 24992 17306 25056
rect 16910 24991 17306 24992
rect 22910 25056 23306 25057
rect 22910 24992 22916 25056
rect 22980 24992 22996 25056
rect 23060 24992 23076 25056
rect 23140 24992 23156 25056
rect 23220 24992 23236 25056
rect 23300 24992 23306 25056
rect 22910 24991 23306 24992
rect 28910 25056 29306 25057
rect 28910 24992 28916 25056
rect 28980 24992 28996 25056
rect 29060 24992 29076 25056
rect 29140 24992 29156 25056
rect 29220 24992 29236 25056
rect 29300 24992 29306 25056
rect 28910 24991 29306 24992
rect 10685 24714 10751 24717
rect 31109 24714 31175 24717
rect 10685 24712 31175 24714
rect 10685 24656 10690 24712
rect 10746 24656 31114 24712
rect 31170 24656 31175 24712
rect 10685 24654 31175 24656
rect 10685 24651 10751 24654
rect 31109 24651 31175 24654
rect 0 24578 800 24608
rect 933 24578 999 24581
rect 0 24576 999 24578
rect 0 24520 938 24576
rect 994 24520 999 24576
rect 0 24518 999 24520
rect 0 24488 800 24518
rect 933 24515 999 24518
rect 4170 24512 4566 24513
rect 4170 24448 4176 24512
rect 4240 24448 4256 24512
rect 4320 24448 4336 24512
rect 4400 24448 4416 24512
rect 4480 24448 4496 24512
rect 4560 24448 4566 24512
rect 4170 24447 4566 24448
rect 10170 24512 10566 24513
rect 10170 24448 10176 24512
rect 10240 24448 10256 24512
rect 10320 24448 10336 24512
rect 10400 24448 10416 24512
rect 10480 24448 10496 24512
rect 10560 24448 10566 24512
rect 10170 24447 10566 24448
rect 16170 24512 16566 24513
rect 16170 24448 16176 24512
rect 16240 24448 16256 24512
rect 16320 24448 16336 24512
rect 16400 24448 16416 24512
rect 16480 24448 16496 24512
rect 16560 24448 16566 24512
rect 16170 24447 16566 24448
rect 22170 24512 22566 24513
rect 22170 24448 22176 24512
rect 22240 24448 22256 24512
rect 22320 24448 22336 24512
rect 22400 24448 22416 24512
rect 22480 24448 22496 24512
rect 22560 24448 22566 24512
rect 22170 24447 22566 24448
rect 28170 24512 28566 24513
rect 28170 24448 28176 24512
rect 28240 24448 28256 24512
rect 28320 24448 28336 24512
rect 28400 24448 28416 24512
rect 28480 24448 28496 24512
rect 28560 24448 28566 24512
rect 28170 24447 28566 24448
rect 4910 23968 5306 23969
rect 4910 23904 4916 23968
rect 4980 23904 4996 23968
rect 5060 23904 5076 23968
rect 5140 23904 5156 23968
rect 5220 23904 5236 23968
rect 5300 23904 5306 23968
rect 4910 23903 5306 23904
rect 10910 23968 11306 23969
rect 10910 23904 10916 23968
rect 10980 23904 10996 23968
rect 11060 23904 11076 23968
rect 11140 23904 11156 23968
rect 11220 23904 11236 23968
rect 11300 23904 11306 23968
rect 10910 23903 11306 23904
rect 16910 23968 17306 23969
rect 16910 23904 16916 23968
rect 16980 23904 16996 23968
rect 17060 23904 17076 23968
rect 17140 23904 17156 23968
rect 17220 23904 17236 23968
rect 17300 23904 17306 23968
rect 16910 23903 17306 23904
rect 22910 23968 23306 23969
rect 22910 23904 22916 23968
rect 22980 23904 22996 23968
rect 23060 23904 23076 23968
rect 23140 23904 23156 23968
rect 23220 23904 23236 23968
rect 23300 23904 23306 23968
rect 22910 23903 23306 23904
rect 28910 23968 29306 23969
rect 28910 23904 28916 23968
rect 28980 23904 28996 23968
rect 29060 23904 29076 23968
rect 29140 23904 29156 23968
rect 29220 23904 29236 23968
rect 29300 23904 29306 23968
rect 28910 23903 29306 23904
rect 14089 23490 14155 23493
rect 14222 23490 14228 23492
rect 14089 23488 14228 23490
rect 14089 23432 14094 23488
rect 14150 23432 14228 23488
rect 14089 23430 14228 23432
rect 14089 23427 14155 23430
rect 14222 23428 14228 23430
rect 14292 23428 14298 23492
rect 4170 23424 4566 23425
rect 4170 23360 4176 23424
rect 4240 23360 4256 23424
rect 4320 23360 4336 23424
rect 4400 23360 4416 23424
rect 4480 23360 4496 23424
rect 4560 23360 4566 23424
rect 4170 23359 4566 23360
rect 10170 23424 10566 23425
rect 10170 23360 10176 23424
rect 10240 23360 10256 23424
rect 10320 23360 10336 23424
rect 10400 23360 10416 23424
rect 10480 23360 10496 23424
rect 10560 23360 10566 23424
rect 10170 23359 10566 23360
rect 16170 23424 16566 23425
rect 16170 23360 16176 23424
rect 16240 23360 16256 23424
rect 16320 23360 16336 23424
rect 16400 23360 16416 23424
rect 16480 23360 16496 23424
rect 16560 23360 16566 23424
rect 16170 23359 16566 23360
rect 22170 23424 22566 23425
rect 22170 23360 22176 23424
rect 22240 23360 22256 23424
rect 22320 23360 22336 23424
rect 22400 23360 22416 23424
rect 22480 23360 22496 23424
rect 22560 23360 22566 23424
rect 22170 23359 22566 23360
rect 28170 23424 28566 23425
rect 28170 23360 28176 23424
rect 28240 23360 28256 23424
rect 28320 23360 28336 23424
rect 28400 23360 28416 23424
rect 28480 23360 28496 23424
rect 28560 23360 28566 23424
rect 28170 23359 28566 23360
rect 4910 22880 5306 22881
rect 4910 22816 4916 22880
rect 4980 22816 4996 22880
rect 5060 22816 5076 22880
rect 5140 22816 5156 22880
rect 5220 22816 5236 22880
rect 5300 22816 5306 22880
rect 4910 22815 5306 22816
rect 10910 22880 11306 22881
rect 10910 22816 10916 22880
rect 10980 22816 10996 22880
rect 11060 22816 11076 22880
rect 11140 22816 11156 22880
rect 11220 22816 11236 22880
rect 11300 22816 11306 22880
rect 10910 22815 11306 22816
rect 16910 22880 17306 22881
rect 16910 22816 16916 22880
rect 16980 22816 16996 22880
rect 17060 22816 17076 22880
rect 17140 22816 17156 22880
rect 17220 22816 17236 22880
rect 17300 22816 17306 22880
rect 16910 22815 17306 22816
rect 22910 22880 23306 22881
rect 22910 22816 22916 22880
rect 22980 22816 22996 22880
rect 23060 22816 23076 22880
rect 23140 22816 23156 22880
rect 23220 22816 23236 22880
rect 23300 22816 23306 22880
rect 22910 22815 23306 22816
rect 28910 22880 29306 22881
rect 28910 22816 28916 22880
rect 28980 22816 28996 22880
rect 29060 22816 29076 22880
rect 29140 22816 29156 22880
rect 29220 22816 29236 22880
rect 29300 22816 29306 22880
rect 28910 22815 29306 22816
rect 4170 22336 4566 22337
rect 4170 22272 4176 22336
rect 4240 22272 4256 22336
rect 4320 22272 4336 22336
rect 4400 22272 4416 22336
rect 4480 22272 4496 22336
rect 4560 22272 4566 22336
rect 4170 22271 4566 22272
rect 10170 22336 10566 22337
rect 10170 22272 10176 22336
rect 10240 22272 10256 22336
rect 10320 22272 10336 22336
rect 10400 22272 10416 22336
rect 10480 22272 10496 22336
rect 10560 22272 10566 22336
rect 10170 22271 10566 22272
rect 16170 22336 16566 22337
rect 16170 22272 16176 22336
rect 16240 22272 16256 22336
rect 16320 22272 16336 22336
rect 16400 22272 16416 22336
rect 16480 22272 16496 22336
rect 16560 22272 16566 22336
rect 16170 22271 16566 22272
rect 22170 22336 22566 22337
rect 22170 22272 22176 22336
rect 22240 22272 22256 22336
rect 22320 22272 22336 22336
rect 22400 22272 22416 22336
rect 22480 22272 22496 22336
rect 22560 22272 22566 22336
rect 22170 22271 22566 22272
rect 28170 22336 28566 22337
rect 28170 22272 28176 22336
rect 28240 22272 28256 22336
rect 28320 22272 28336 22336
rect 28400 22272 28416 22336
rect 28480 22272 28496 22336
rect 28560 22272 28566 22336
rect 28170 22271 28566 22272
rect 4910 21792 5306 21793
rect 4910 21728 4916 21792
rect 4980 21728 4996 21792
rect 5060 21728 5076 21792
rect 5140 21728 5156 21792
rect 5220 21728 5236 21792
rect 5300 21728 5306 21792
rect 4910 21727 5306 21728
rect 10910 21792 11306 21793
rect 10910 21728 10916 21792
rect 10980 21728 10996 21792
rect 11060 21728 11076 21792
rect 11140 21728 11156 21792
rect 11220 21728 11236 21792
rect 11300 21728 11306 21792
rect 10910 21727 11306 21728
rect 16910 21792 17306 21793
rect 16910 21728 16916 21792
rect 16980 21728 16996 21792
rect 17060 21728 17076 21792
rect 17140 21728 17156 21792
rect 17220 21728 17236 21792
rect 17300 21728 17306 21792
rect 16910 21727 17306 21728
rect 22910 21792 23306 21793
rect 22910 21728 22916 21792
rect 22980 21728 22996 21792
rect 23060 21728 23076 21792
rect 23140 21728 23156 21792
rect 23220 21728 23236 21792
rect 23300 21728 23306 21792
rect 22910 21727 23306 21728
rect 28910 21792 29306 21793
rect 28910 21728 28916 21792
rect 28980 21728 28996 21792
rect 29060 21728 29076 21792
rect 29140 21728 29156 21792
rect 29220 21728 29236 21792
rect 29300 21728 29306 21792
rect 28910 21727 29306 21728
rect 8201 21586 8267 21589
rect 11329 21586 11395 21589
rect 8201 21584 11395 21586
rect 8201 21528 8206 21584
rect 8262 21528 11334 21584
rect 11390 21528 11395 21584
rect 8201 21526 11395 21528
rect 8201 21523 8267 21526
rect 11329 21523 11395 21526
rect 20713 21586 20779 21589
rect 24853 21586 24919 21589
rect 20713 21584 24919 21586
rect 20713 21528 20718 21584
rect 20774 21528 24858 21584
rect 24914 21528 24919 21584
rect 20713 21526 24919 21528
rect 20713 21523 20779 21526
rect 24853 21523 24919 21526
rect 4170 21248 4566 21249
rect 4170 21184 4176 21248
rect 4240 21184 4256 21248
rect 4320 21184 4336 21248
rect 4400 21184 4416 21248
rect 4480 21184 4496 21248
rect 4560 21184 4566 21248
rect 4170 21183 4566 21184
rect 10170 21248 10566 21249
rect 10170 21184 10176 21248
rect 10240 21184 10256 21248
rect 10320 21184 10336 21248
rect 10400 21184 10416 21248
rect 10480 21184 10496 21248
rect 10560 21184 10566 21248
rect 10170 21183 10566 21184
rect 16170 21248 16566 21249
rect 16170 21184 16176 21248
rect 16240 21184 16256 21248
rect 16320 21184 16336 21248
rect 16400 21184 16416 21248
rect 16480 21184 16496 21248
rect 16560 21184 16566 21248
rect 16170 21183 16566 21184
rect 22170 21248 22566 21249
rect 22170 21184 22176 21248
rect 22240 21184 22256 21248
rect 22320 21184 22336 21248
rect 22400 21184 22416 21248
rect 22480 21184 22496 21248
rect 22560 21184 22566 21248
rect 22170 21183 22566 21184
rect 28170 21248 28566 21249
rect 28170 21184 28176 21248
rect 28240 21184 28256 21248
rect 28320 21184 28336 21248
rect 28400 21184 28416 21248
rect 28480 21184 28496 21248
rect 28560 21184 28566 21248
rect 28170 21183 28566 21184
rect 12157 20770 12223 20773
rect 20713 20772 20779 20773
rect 12934 20770 12940 20772
rect 12157 20768 12940 20770
rect 12157 20712 12162 20768
rect 12218 20712 12940 20768
rect 12157 20710 12940 20712
rect 12157 20707 12223 20710
rect 12934 20708 12940 20710
rect 13004 20708 13010 20772
rect 20662 20708 20668 20772
rect 20732 20770 20779 20772
rect 20732 20768 20824 20770
rect 20774 20712 20824 20768
rect 20732 20710 20824 20712
rect 20732 20708 20779 20710
rect 20713 20707 20779 20708
rect 4910 20704 5306 20705
rect 4910 20640 4916 20704
rect 4980 20640 4996 20704
rect 5060 20640 5076 20704
rect 5140 20640 5156 20704
rect 5220 20640 5236 20704
rect 5300 20640 5306 20704
rect 4910 20639 5306 20640
rect 10910 20704 11306 20705
rect 10910 20640 10916 20704
rect 10980 20640 10996 20704
rect 11060 20640 11076 20704
rect 11140 20640 11156 20704
rect 11220 20640 11236 20704
rect 11300 20640 11306 20704
rect 10910 20639 11306 20640
rect 16910 20704 17306 20705
rect 16910 20640 16916 20704
rect 16980 20640 16996 20704
rect 17060 20640 17076 20704
rect 17140 20640 17156 20704
rect 17220 20640 17236 20704
rect 17300 20640 17306 20704
rect 16910 20639 17306 20640
rect 22910 20704 23306 20705
rect 22910 20640 22916 20704
rect 22980 20640 22996 20704
rect 23060 20640 23076 20704
rect 23140 20640 23156 20704
rect 23220 20640 23236 20704
rect 23300 20640 23306 20704
rect 22910 20639 23306 20640
rect 28910 20704 29306 20705
rect 28910 20640 28916 20704
rect 28980 20640 28996 20704
rect 29060 20640 29076 20704
rect 29140 20640 29156 20704
rect 29220 20640 29236 20704
rect 29300 20640 29306 20704
rect 28910 20639 29306 20640
rect 4170 20160 4566 20161
rect 4170 20096 4176 20160
rect 4240 20096 4256 20160
rect 4320 20096 4336 20160
rect 4400 20096 4416 20160
rect 4480 20096 4496 20160
rect 4560 20096 4566 20160
rect 4170 20095 4566 20096
rect 10170 20160 10566 20161
rect 10170 20096 10176 20160
rect 10240 20096 10256 20160
rect 10320 20096 10336 20160
rect 10400 20096 10416 20160
rect 10480 20096 10496 20160
rect 10560 20096 10566 20160
rect 10170 20095 10566 20096
rect 16170 20160 16566 20161
rect 16170 20096 16176 20160
rect 16240 20096 16256 20160
rect 16320 20096 16336 20160
rect 16400 20096 16416 20160
rect 16480 20096 16496 20160
rect 16560 20096 16566 20160
rect 16170 20095 16566 20096
rect 22170 20160 22566 20161
rect 22170 20096 22176 20160
rect 22240 20096 22256 20160
rect 22320 20096 22336 20160
rect 22400 20096 22416 20160
rect 22480 20096 22496 20160
rect 22560 20096 22566 20160
rect 22170 20095 22566 20096
rect 28170 20160 28566 20161
rect 28170 20096 28176 20160
rect 28240 20096 28256 20160
rect 28320 20096 28336 20160
rect 28400 20096 28416 20160
rect 28480 20096 28496 20160
rect 28560 20096 28566 20160
rect 28170 20095 28566 20096
rect 31845 19818 31911 19821
rect 32174 19818 32974 19848
rect 31845 19816 32974 19818
rect 31845 19760 31850 19816
rect 31906 19760 32974 19816
rect 31845 19758 32974 19760
rect 31845 19755 31911 19758
rect 32174 19728 32974 19758
rect 4910 19616 5306 19617
rect 4910 19552 4916 19616
rect 4980 19552 4996 19616
rect 5060 19552 5076 19616
rect 5140 19552 5156 19616
rect 5220 19552 5236 19616
rect 5300 19552 5306 19616
rect 4910 19551 5306 19552
rect 10910 19616 11306 19617
rect 10910 19552 10916 19616
rect 10980 19552 10996 19616
rect 11060 19552 11076 19616
rect 11140 19552 11156 19616
rect 11220 19552 11236 19616
rect 11300 19552 11306 19616
rect 10910 19551 11306 19552
rect 16910 19616 17306 19617
rect 16910 19552 16916 19616
rect 16980 19552 16996 19616
rect 17060 19552 17076 19616
rect 17140 19552 17156 19616
rect 17220 19552 17236 19616
rect 17300 19552 17306 19616
rect 16910 19551 17306 19552
rect 22910 19616 23306 19617
rect 22910 19552 22916 19616
rect 22980 19552 22996 19616
rect 23060 19552 23076 19616
rect 23140 19552 23156 19616
rect 23220 19552 23236 19616
rect 23300 19552 23306 19616
rect 22910 19551 23306 19552
rect 28910 19616 29306 19617
rect 28910 19552 28916 19616
rect 28980 19552 28996 19616
rect 29060 19552 29076 19616
rect 29140 19552 29156 19616
rect 29220 19552 29236 19616
rect 29300 19552 29306 19616
rect 28910 19551 29306 19552
rect 14222 19348 14228 19412
rect 14292 19410 14298 19412
rect 14365 19410 14431 19413
rect 14292 19408 14431 19410
rect 14292 19352 14370 19408
rect 14426 19352 14431 19408
rect 14292 19350 14431 19352
rect 14292 19348 14298 19350
rect 14365 19347 14431 19350
rect 4170 19072 4566 19073
rect 4170 19008 4176 19072
rect 4240 19008 4256 19072
rect 4320 19008 4336 19072
rect 4400 19008 4416 19072
rect 4480 19008 4496 19072
rect 4560 19008 4566 19072
rect 4170 19007 4566 19008
rect 10170 19072 10566 19073
rect 10170 19008 10176 19072
rect 10240 19008 10256 19072
rect 10320 19008 10336 19072
rect 10400 19008 10416 19072
rect 10480 19008 10496 19072
rect 10560 19008 10566 19072
rect 10170 19007 10566 19008
rect 16170 19072 16566 19073
rect 16170 19008 16176 19072
rect 16240 19008 16256 19072
rect 16320 19008 16336 19072
rect 16400 19008 16416 19072
rect 16480 19008 16496 19072
rect 16560 19008 16566 19072
rect 16170 19007 16566 19008
rect 22170 19072 22566 19073
rect 22170 19008 22176 19072
rect 22240 19008 22256 19072
rect 22320 19008 22336 19072
rect 22400 19008 22416 19072
rect 22480 19008 22496 19072
rect 22560 19008 22566 19072
rect 22170 19007 22566 19008
rect 28170 19072 28566 19073
rect 28170 19008 28176 19072
rect 28240 19008 28256 19072
rect 28320 19008 28336 19072
rect 28400 19008 28416 19072
rect 28480 19008 28496 19072
rect 28560 19008 28566 19072
rect 28170 19007 28566 19008
rect 4910 18528 5306 18529
rect 0 18458 800 18488
rect 4910 18464 4916 18528
rect 4980 18464 4996 18528
rect 5060 18464 5076 18528
rect 5140 18464 5156 18528
rect 5220 18464 5236 18528
rect 5300 18464 5306 18528
rect 4910 18463 5306 18464
rect 10910 18528 11306 18529
rect 10910 18464 10916 18528
rect 10980 18464 10996 18528
rect 11060 18464 11076 18528
rect 11140 18464 11156 18528
rect 11220 18464 11236 18528
rect 11300 18464 11306 18528
rect 10910 18463 11306 18464
rect 16910 18528 17306 18529
rect 16910 18464 16916 18528
rect 16980 18464 16996 18528
rect 17060 18464 17076 18528
rect 17140 18464 17156 18528
rect 17220 18464 17236 18528
rect 17300 18464 17306 18528
rect 16910 18463 17306 18464
rect 22910 18528 23306 18529
rect 22910 18464 22916 18528
rect 22980 18464 22996 18528
rect 23060 18464 23076 18528
rect 23140 18464 23156 18528
rect 23220 18464 23236 18528
rect 23300 18464 23306 18528
rect 22910 18463 23306 18464
rect 28910 18528 29306 18529
rect 28910 18464 28916 18528
rect 28980 18464 28996 18528
rect 29060 18464 29076 18528
rect 29140 18464 29156 18528
rect 29220 18464 29236 18528
rect 29300 18464 29306 18528
rect 28910 18463 29306 18464
rect 933 18458 999 18461
rect 0 18456 999 18458
rect 0 18400 938 18456
rect 994 18400 999 18456
rect 0 18398 999 18400
rect 0 18368 800 18398
rect 933 18395 999 18398
rect 4170 17984 4566 17985
rect 4170 17920 4176 17984
rect 4240 17920 4256 17984
rect 4320 17920 4336 17984
rect 4400 17920 4416 17984
rect 4480 17920 4496 17984
rect 4560 17920 4566 17984
rect 4170 17919 4566 17920
rect 10170 17984 10566 17985
rect 10170 17920 10176 17984
rect 10240 17920 10256 17984
rect 10320 17920 10336 17984
rect 10400 17920 10416 17984
rect 10480 17920 10496 17984
rect 10560 17920 10566 17984
rect 10170 17919 10566 17920
rect 16170 17984 16566 17985
rect 16170 17920 16176 17984
rect 16240 17920 16256 17984
rect 16320 17920 16336 17984
rect 16400 17920 16416 17984
rect 16480 17920 16496 17984
rect 16560 17920 16566 17984
rect 16170 17919 16566 17920
rect 22170 17984 22566 17985
rect 22170 17920 22176 17984
rect 22240 17920 22256 17984
rect 22320 17920 22336 17984
rect 22400 17920 22416 17984
rect 22480 17920 22496 17984
rect 22560 17920 22566 17984
rect 22170 17919 22566 17920
rect 28170 17984 28566 17985
rect 28170 17920 28176 17984
rect 28240 17920 28256 17984
rect 28320 17920 28336 17984
rect 28400 17920 28416 17984
rect 28480 17920 28496 17984
rect 28560 17920 28566 17984
rect 28170 17919 28566 17920
rect 18413 17642 18479 17645
rect 27838 17642 27844 17644
rect 18413 17640 27844 17642
rect 18413 17584 18418 17640
rect 18474 17584 27844 17640
rect 18413 17582 27844 17584
rect 18413 17579 18479 17582
rect 27838 17580 27844 17582
rect 27908 17580 27914 17644
rect 17861 17506 17927 17509
rect 19374 17506 19380 17508
rect 17861 17504 19380 17506
rect 17861 17448 17866 17504
rect 17922 17448 19380 17504
rect 17861 17446 19380 17448
rect 17861 17443 17927 17446
rect 19374 17444 19380 17446
rect 19444 17506 19450 17508
rect 20662 17506 20668 17508
rect 19444 17446 20668 17506
rect 19444 17444 19450 17446
rect 20662 17444 20668 17446
rect 20732 17444 20738 17508
rect 4910 17440 5306 17441
rect 4910 17376 4916 17440
rect 4980 17376 4996 17440
rect 5060 17376 5076 17440
rect 5140 17376 5156 17440
rect 5220 17376 5236 17440
rect 5300 17376 5306 17440
rect 4910 17375 5306 17376
rect 10910 17440 11306 17441
rect 10910 17376 10916 17440
rect 10980 17376 10996 17440
rect 11060 17376 11076 17440
rect 11140 17376 11156 17440
rect 11220 17376 11236 17440
rect 11300 17376 11306 17440
rect 10910 17375 11306 17376
rect 16910 17440 17306 17441
rect 16910 17376 16916 17440
rect 16980 17376 16996 17440
rect 17060 17376 17076 17440
rect 17140 17376 17156 17440
rect 17220 17376 17236 17440
rect 17300 17376 17306 17440
rect 16910 17375 17306 17376
rect 22910 17440 23306 17441
rect 22910 17376 22916 17440
rect 22980 17376 22996 17440
rect 23060 17376 23076 17440
rect 23140 17376 23156 17440
rect 23220 17376 23236 17440
rect 23300 17376 23306 17440
rect 22910 17375 23306 17376
rect 28910 17440 29306 17441
rect 28910 17376 28916 17440
rect 28980 17376 28996 17440
rect 29060 17376 29076 17440
rect 29140 17376 29156 17440
rect 29220 17376 29236 17440
rect 29300 17376 29306 17440
rect 28910 17375 29306 17376
rect 4170 16896 4566 16897
rect 4170 16832 4176 16896
rect 4240 16832 4256 16896
rect 4320 16832 4336 16896
rect 4400 16832 4416 16896
rect 4480 16832 4496 16896
rect 4560 16832 4566 16896
rect 4170 16831 4566 16832
rect 10170 16896 10566 16897
rect 10170 16832 10176 16896
rect 10240 16832 10256 16896
rect 10320 16832 10336 16896
rect 10400 16832 10416 16896
rect 10480 16832 10496 16896
rect 10560 16832 10566 16896
rect 10170 16831 10566 16832
rect 16170 16896 16566 16897
rect 16170 16832 16176 16896
rect 16240 16832 16256 16896
rect 16320 16832 16336 16896
rect 16400 16832 16416 16896
rect 16480 16832 16496 16896
rect 16560 16832 16566 16896
rect 16170 16831 16566 16832
rect 22170 16896 22566 16897
rect 22170 16832 22176 16896
rect 22240 16832 22256 16896
rect 22320 16832 22336 16896
rect 22400 16832 22416 16896
rect 22480 16832 22496 16896
rect 22560 16832 22566 16896
rect 22170 16831 22566 16832
rect 28170 16896 28566 16897
rect 28170 16832 28176 16896
rect 28240 16832 28256 16896
rect 28320 16832 28336 16896
rect 28400 16832 28416 16896
rect 28480 16832 28496 16896
rect 28560 16832 28566 16896
rect 28170 16831 28566 16832
rect 29085 16690 29151 16693
rect 30925 16690 30991 16693
rect 29085 16688 30991 16690
rect 29085 16632 29090 16688
rect 29146 16632 30930 16688
rect 30986 16632 30991 16688
rect 29085 16630 30991 16632
rect 29085 16627 29151 16630
rect 30925 16627 30991 16630
rect 4910 16352 5306 16353
rect 4910 16288 4916 16352
rect 4980 16288 4996 16352
rect 5060 16288 5076 16352
rect 5140 16288 5156 16352
rect 5220 16288 5236 16352
rect 5300 16288 5306 16352
rect 4910 16287 5306 16288
rect 10910 16352 11306 16353
rect 10910 16288 10916 16352
rect 10980 16288 10996 16352
rect 11060 16288 11076 16352
rect 11140 16288 11156 16352
rect 11220 16288 11236 16352
rect 11300 16288 11306 16352
rect 10910 16287 11306 16288
rect 16910 16352 17306 16353
rect 16910 16288 16916 16352
rect 16980 16288 16996 16352
rect 17060 16288 17076 16352
rect 17140 16288 17156 16352
rect 17220 16288 17236 16352
rect 17300 16288 17306 16352
rect 16910 16287 17306 16288
rect 22910 16352 23306 16353
rect 22910 16288 22916 16352
rect 22980 16288 22996 16352
rect 23060 16288 23076 16352
rect 23140 16288 23156 16352
rect 23220 16288 23236 16352
rect 23300 16288 23306 16352
rect 22910 16287 23306 16288
rect 28910 16352 29306 16353
rect 28910 16288 28916 16352
rect 28980 16288 28996 16352
rect 29060 16288 29076 16352
rect 29140 16288 29156 16352
rect 29220 16288 29236 16352
rect 29300 16288 29306 16352
rect 28910 16287 29306 16288
rect 21357 16010 21423 16013
rect 22921 16010 22987 16013
rect 23841 16010 23907 16013
rect 21357 16008 23907 16010
rect 21357 15952 21362 16008
rect 21418 15952 22926 16008
rect 22982 15952 23846 16008
rect 23902 15952 23907 16008
rect 21357 15950 23907 15952
rect 21357 15947 21423 15950
rect 22921 15947 22987 15950
rect 23841 15947 23907 15950
rect 4170 15808 4566 15809
rect 4170 15744 4176 15808
rect 4240 15744 4256 15808
rect 4320 15744 4336 15808
rect 4400 15744 4416 15808
rect 4480 15744 4496 15808
rect 4560 15744 4566 15808
rect 4170 15743 4566 15744
rect 10170 15808 10566 15809
rect 10170 15744 10176 15808
rect 10240 15744 10256 15808
rect 10320 15744 10336 15808
rect 10400 15744 10416 15808
rect 10480 15744 10496 15808
rect 10560 15744 10566 15808
rect 10170 15743 10566 15744
rect 16170 15808 16566 15809
rect 16170 15744 16176 15808
rect 16240 15744 16256 15808
rect 16320 15744 16336 15808
rect 16400 15744 16416 15808
rect 16480 15744 16496 15808
rect 16560 15744 16566 15808
rect 16170 15743 16566 15744
rect 22170 15808 22566 15809
rect 22170 15744 22176 15808
rect 22240 15744 22256 15808
rect 22320 15744 22336 15808
rect 22400 15744 22416 15808
rect 22480 15744 22496 15808
rect 22560 15744 22566 15808
rect 22170 15743 22566 15744
rect 28170 15808 28566 15809
rect 28170 15744 28176 15808
rect 28240 15744 28256 15808
rect 28320 15744 28336 15808
rect 28400 15744 28416 15808
rect 28480 15744 28496 15808
rect 28560 15744 28566 15808
rect 28170 15743 28566 15744
rect 4910 15264 5306 15265
rect 4910 15200 4916 15264
rect 4980 15200 4996 15264
rect 5060 15200 5076 15264
rect 5140 15200 5156 15264
rect 5220 15200 5236 15264
rect 5300 15200 5306 15264
rect 4910 15199 5306 15200
rect 10910 15264 11306 15265
rect 10910 15200 10916 15264
rect 10980 15200 10996 15264
rect 11060 15200 11076 15264
rect 11140 15200 11156 15264
rect 11220 15200 11236 15264
rect 11300 15200 11306 15264
rect 10910 15199 11306 15200
rect 16910 15264 17306 15265
rect 16910 15200 16916 15264
rect 16980 15200 16996 15264
rect 17060 15200 17076 15264
rect 17140 15200 17156 15264
rect 17220 15200 17236 15264
rect 17300 15200 17306 15264
rect 16910 15199 17306 15200
rect 22910 15264 23306 15265
rect 22910 15200 22916 15264
rect 22980 15200 22996 15264
rect 23060 15200 23076 15264
rect 23140 15200 23156 15264
rect 23220 15200 23236 15264
rect 23300 15200 23306 15264
rect 22910 15199 23306 15200
rect 28910 15264 29306 15265
rect 28910 15200 28916 15264
rect 28980 15200 28996 15264
rect 29060 15200 29076 15264
rect 29140 15200 29156 15264
rect 29220 15200 29236 15264
rect 29300 15200 29306 15264
rect 28910 15199 29306 15200
rect 4170 14720 4566 14721
rect 4170 14656 4176 14720
rect 4240 14656 4256 14720
rect 4320 14656 4336 14720
rect 4400 14656 4416 14720
rect 4480 14656 4496 14720
rect 4560 14656 4566 14720
rect 4170 14655 4566 14656
rect 10170 14720 10566 14721
rect 10170 14656 10176 14720
rect 10240 14656 10256 14720
rect 10320 14656 10336 14720
rect 10400 14656 10416 14720
rect 10480 14656 10496 14720
rect 10560 14656 10566 14720
rect 10170 14655 10566 14656
rect 16170 14720 16566 14721
rect 16170 14656 16176 14720
rect 16240 14656 16256 14720
rect 16320 14656 16336 14720
rect 16400 14656 16416 14720
rect 16480 14656 16496 14720
rect 16560 14656 16566 14720
rect 16170 14655 16566 14656
rect 22170 14720 22566 14721
rect 22170 14656 22176 14720
rect 22240 14656 22256 14720
rect 22320 14656 22336 14720
rect 22400 14656 22416 14720
rect 22480 14656 22496 14720
rect 22560 14656 22566 14720
rect 22170 14655 22566 14656
rect 28170 14720 28566 14721
rect 28170 14656 28176 14720
rect 28240 14656 28256 14720
rect 28320 14656 28336 14720
rect 28400 14656 28416 14720
rect 28480 14656 28496 14720
rect 28560 14656 28566 14720
rect 28170 14655 28566 14656
rect 4910 14176 5306 14177
rect 4910 14112 4916 14176
rect 4980 14112 4996 14176
rect 5060 14112 5076 14176
rect 5140 14112 5156 14176
rect 5220 14112 5236 14176
rect 5300 14112 5306 14176
rect 4910 14111 5306 14112
rect 10910 14176 11306 14177
rect 10910 14112 10916 14176
rect 10980 14112 10996 14176
rect 11060 14112 11076 14176
rect 11140 14112 11156 14176
rect 11220 14112 11236 14176
rect 11300 14112 11306 14176
rect 10910 14111 11306 14112
rect 16910 14176 17306 14177
rect 16910 14112 16916 14176
rect 16980 14112 16996 14176
rect 17060 14112 17076 14176
rect 17140 14112 17156 14176
rect 17220 14112 17236 14176
rect 17300 14112 17306 14176
rect 16910 14111 17306 14112
rect 22910 14176 23306 14177
rect 22910 14112 22916 14176
rect 22980 14112 22996 14176
rect 23060 14112 23076 14176
rect 23140 14112 23156 14176
rect 23220 14112 23236 14176
rect 23300 14112 23306 14176
rect 22910 14111 23306 14112
rect 28910 14176 29306 14177
rect 28910 14112 28916 14176
rect 28980 14112 28996 14176
rect 29060 14112 29076 14176
rect 29140 14112 29156 14176
rect 29220 14112 29236 14176
rect 29300 14112 29306 14176
rect 28910 14111 29306 14112
rect 31477 13698 31543 13701
rect 32174 13698 32974 13728
rect 31477 13696 32974 13698
rect 31477 13640 31482 13696
rect 31538 13640 32974 13696
rect 31477 13638 32974 13640
rect 31477 13635 31543 13638
rect 4170 13632 4566 13633
rect 4170 13568 4176 13632
rect 4240 13568 4256 13632
rect 4320 13568 4336 13632
rect 4400 13568 4416 13632
rect 4480 13568 4496 13632
rect 4560 13568 4566 13632
rect 4170 13567 4566 13568
rect 10170 13632 10566 13633
rect 10170 13568 10176 13632
rect 10240 13568 10256 13632
rect 10320 13568 10336 13632
rect 10400 13568 10416 13632
rect 10480 13568 10496 13632
rect 10560 13568 10566 13632
rect 10170 13567 10566 13568
rect 16170 13632 16566 13633
rect 16170 13568 16176 13632
rect 16240 13568 16256 13632
rect 16320 13568 16336 13632
rect 16400 13568 16416 13632
rect 16480 13568 16496 13632
rect 16560 13568 16566 13632
rect 16170 13567 16566 13568
rect 22170 13632 22566 13633
rect 22170 13568 22176 13632
rect 22240 13568 22256 13632
rect 22320 13568 22336 13632
rect 22400 13568 22416 13632
rect 22480 13568 22496 13632
rect 22560 13568 22566 13632
rect 22170 13567 22566 13568
rect 28170 13632 28566 13633
rect 28170 13568 28176 13632
rect 28240 13568 28256 13632
rect 28320 13568 28336 13632
rect 28400 13568 28416 13632
rect 28480 13568 28496 13632
rect 28560 13568 28566 13632
rect 32174 13608 32974 13638
rect 28170 13567 28566 13568
rect 4910 13088 5306 13089
rect 4910 13024 4916 13088
rect 4980 13024 4996 13088
rect 5060 13024 5076 13088
rect 5140 13024 5156 13088
rect 5220 13024 5236 13088
rect 5300 13024 5306 13088
rect 4910 13023 5306 13024
rect 10910 13088 11306 13089
rect 10910 13024 10916 13088
rect 10980 13024 10996 13088
rect 11060 13024 11076 13088
rect 11140 13024 11156 13088
rect 11220 13024 11236 13088
rect 11300 13024 11306 13088
rect 10910 13023 11306 13024
rect 16910 13088 17306 13089
rect 16910 13024 16916 13088
rect 16980 13024 16996 13088
rect 17060 13024 17076 13088
rect 17140 13024 17156 13088
rect 17220 13024 17236 13088
rect 17300 13024 17306 13088
rect 16910 13023 17306 13024
rect 22910 13088 23306 13089
rect 22910 13024 22916 13088
rect 22980 13024 22996 13088
rect 23060 13024 23076 13088
rect 23140 13024 23156 13088
rect 23220 13024 23236 13088
rect 23300 13024 23306 13088
rect 22910 13023 23306 13024
rect 28910 13088 29306 13089
rect 28910 13024 28916 13088
rect 28980 13024 28996 13088
rect 29060 13024 29076 13088
rect 29140 13024 29156 13088
rect 29220 13024 29236 13088
rect 29300 13024 29306 13088
rect 28910 13023 29306 13024
rect 12934 12684 12940 12748
rect 13004 12746 13010 12748
rect 19374 12746 19380 12748
rect 13004 12686 19380 12746
rect 13004 12684 13010 12686
rect 19374 12684 19380 12686
rect 19444 12746 19450 12748
rect 20437 12746 20503 12749
rect 19444 12744 20503 12746
rect 19444 12688 20442 12744
rect 20498 12688 20503 12744
rect 19444 12686 20503 12688
rect 19444 12684 19450 12686
rect 20437 12683 20503 12686
rect 4170 12544 4566 12545
rect 4170 12480 4176 12544
rect 4240 12480 4256 12544
rect 4320 12480 4336 12544
rect 4400 12480 4416 12544
rect 4480 12480 4496 12544
rect 4560 12480 4566 12544
rect 4170 12479 4566 12480
rect 10170 12544 10566 12545
rect 10170 12480 10176 12544
rect 10240 12480 10256 12544
rect 10320 12480 10336 12544
rect 10400 12480 10416 12544
rect 10480 12480 10496 12544
rect 10560 12480 10566 12544
rect 10170 12479 10566 12480
rect 16170 12544 16566 12545
rect 16170 12480 16176 12544
rect 16240 12480 16256 12544
rect 16320 12480 16336 12544
rect 16400 12480 16416 12544
rect 16480 12480 16496 12544
rect 16560 12480 16566 12544
rect 16170 12479 16566 12480
rect 22170 12544 22566 12545
rect 22170 12480 22176 12544
rect 22240 12480 22256 12544
rect 22320 12480 22336 12544
rect 22400 12480 22416 12544
rect 22480 12480 22496 12544
rect 22560 12480 22566 12544
rect 22170 12479 22566 12480
rect 28170 12544 28566 12545
rect 28170 12480 28176 12544
rect 28240 12480 28256 12544
rect 28320 12480 28336 12544
rect 28400 12480 28416 12544
rect 28480 12480 28496 12544
rect 28560 12480 28566 12544
rect 28170 12479 28566 12480
rect 0 12338 800 12368
rect 1485 12338 1551 12341
rect 0 12336 1551 12338
rect 0 12280 1490 12336
rect 1546 12280 1551 12336
rect 0 12278 1551 12280
rect 0 12248 800 12278
rect 1485 12275 1551 12278
rect 4910 12000 5306 12001
rect 4910 11936 4916 12000
rect 4980 11936 4996 12000
rect 5060 11936 5076 12000
rect 5140 11936 5156 12000
rect 5220 11936 5236 12000
rect 5300 11936 5306 12000
rect 4910 11935 5306 11936
rect 10910 12000 11306 12001
rect 10910 11936 10916 12000
rect 10980 11936 10996 12000
rect 11060 11936 11076 12000
rect 11140 11936 11156 12000
rect 11220 11936 11236 12000
rect 11300 11936 11306 12000
rect 10910 11935 11306 11936
rect 16910 12000 17306 12001
rect 16910 11936 16916 12000
rect 16980 11936 16996 12000
rect 17060 11936 17076 12000
rect 17140 11936 17156 12000
rect 17220 11936 17236 12000
rect 17300 11936 17306 12000
rect 16910 11935 17306 11936
rect 22910 12000 23306 12001
rect 22910 11936 22916 12000
rect 22980 11936 22996 12000
rect 23060 11936 23076 12000
rect 23140 11936 23156 12000
rect 23220 11936 23236 12000
rect 23300 11936 23306 12000
rect 22910 11935 23306 11936
rect 28910 12000 29306 12001
rect 28910 11936 28916 12000
rect 28980 11936 28996 12000
rect 29060 11936 29076 12000
rect 29140 11936 29156 12000
rect 29220 11936 29236 12000
rect 29300 11936 29306 12000
rect 28910 11935 29306 11936
rect 21633 11794 21699 11797
rect 25405 11794 25471 11797
rect 21633 11792 25471 11794
rect 21633 11736 21638 11792
rect 21694 11736 25410 11792
rect 25466 11736 25471 11792
rect 21633 11734 25471 11736
rect 21633 11731 21699 11734
rect 25405 11731 25471 11734
rect 4170 11456 4566 11457
rect 4170 11392 4176 11456
rect 4240 11392 4256 11456
rect 4320 11392 4336 11456
rect 4400 11392 4416 11456
rect 4480 11392 4496 11456
rect 4560 11392 4566 11456
rect 4170 11391 4566 11392
rect 10170 11456 10566 11457
rect 10170 11392 10176 11456
rect 10240 11392 10256 11456
rect 10320 11392 10336 11456
rect 10400 11392 10416 11456
rect 10480 11392 10496 11456
rect 10560 11392 10566 11456
rect 10170 11391 10566 11392
rect 16170 11456 16566 11457
rect 16170 11392 16176 11456
rect 16240 11392 16256 11456
rect 16320 11392 16336 11456
rect 16400 11392 16416 11456
rect 16480 11392 16496 11456
rect 16560 11392 16566 11456
rect 16170 11391 16566 11392
rect 22170 11456 22566 11457
rect 22170 11392 22176 11456
rect 22240 11392 22256 11456
rect 22320 11392 22336 11456
rect 22400 11392 22416 11456
rect 22480 11392 22496 11456
rect 22560 11392 22566 11456
rect 22170 11391 22566 11392
rect 28170 11456 28566 11457
rect 28170 11392 28176 11456
rect 28240 11392 28256 11456
rect 28320 11392 28336 11456
rect 28400 11392 28416 11456
rect 28480 11392 28496 11456
rect 28560 11392 28566 11456
rect 28170 11391 28566 11392
rect 12985 11388 13051 11389
rect 12934 11324 12940 11388
rect 13004 11386 13051 11388
rect 13004 11384 13096 11386
rect 13046 11328 13096 11384
rect 13004 11326 13096 11328
rect 13004 11324 13051 11326
rect 12985 11323 13051 11324
rect 4910 10912 5306 10913
rect 4910 10848 4916 10912
rect 4980 10848 4996 10912
rect 5060 10848 5076 10912
rect 5140 10848 5156 10912
rect 5220 10848 5236 10912
rect 5300 10848 5306 10912
rect 4910 10847 5306 10848
rect 10910 10912 11306 10913
rect 10910 10848 10916 10912
rect 10980 10848 10996 10912
rect 11060 10848 11076 10912
rect 11140 10848 11156 10912
rect 11220 10848 11236 10912
rect 11300 10848 11306 10912
rect 10910 10847 11306 10848
rect 16910 10912 17306 10913
rect 16910 10848 16916 10912
rect 16980 10848 16996 10912
rect 17060 10848 17076 10912
rect 17140 10848 17156 10912
rect 17220 10848 17236 10912
rect 17300 10848 17306 10912
rect 16910 10847 17306 10848
rect 22910 10912 23306 10913
rect 22910 10848 22916 10912
rect 22980 10848 22996 10912
rect 23060 10848 23076 10912
rect 23140 10848 23156 10912
rect 23220 10848 23236 10912
rect 23300 10848 23306 10912
rect 22910 10847 23306 10848
rect 28910 10912 29306 10913
rect 28910 10848 28916 10912
rect 28980 10848 28996 10912
rect 29060 10848 29076 10912
rect 29140 10848 29156 10912
rect 29220 10848 29236 10912
rect 29300 10848 29306 10912
rect 28910 10847 29306 10848
rect 4170 10368 4566 10369
rect 4170 10304 4176 10368
rect 4240 10304 4256 10368
rect 4320 10304 4336 10368
rect 4400 10304 4416 10368
rect 4480 10304 4496 10368
rect 4560 10304 4566 10368
rect 4170 10303 4566 10304
rect 10170 10368 10566 10369
rect 10170 10304 10176 10368
rect 10240 10304 10256 10368
rect 10320 10304 10336 10368
rect 10400 10304 10416 10368
rect 10480 10304 10496 10368
rect 10560 10304 10566 10368
rect 10170 10303 10566 10304
rect 16170 10368 16566 10369
rect 16170 10304 16176 10368
rect 16240 10304 16256 10368
rect 16320 10304 16336 10368
rect 16400 10304 16416 10368
rect 16480 10304 16496 10368
rect 16560 10304 16566 10368
rect 16170 10303 16566 10304
rect 22170 10368 22566 10369
rect 22170 10304 22176 10368
rect 22240 10304 22256 10368
rect 22320 10304 22336 10368
rect 22400 10304 22416 10368
rect 22480 10304 22496 10368
rect 22560 10304 22566 10368
rect 22170 10303 22566 10304
rect 28170 10368 28566 10369
rect 28170 10304 28176 10368
rect 28240 10304 28256 10368
rect 28320 10304 28336 10368
rect 28400 10304 28416 10368
rect 28480 10304 28496 10368
rect 28560 10304 28566 10368
rect 28170 10303 28566 10304
rect 4910 9824 5306 9825
rect 4910 9760 4916 9824
rect 4980 9760 4996 9824
rect 5060 9760 5076 9824
rect 5140 9760 5156 9824
rect 5220 9760 5236 9824
rect 5300 9760 5306 9824
rect 4910 9759 5306 9760
rect 10910 9824 11306 9825
rect 10910 9760 10916 9824
rect 10980 9760 10996 9824
rect 11060 9760 11076 9824
rect 11140 9760 11156 9824
rect 11220 9760 11236 9824
rect 11300 9760 11306 9824
rect 10910 9759 11306 9760
rect 16910 9824 17306 9825
rect 16910 9760 16916 9824
rect 16980 9760 16996 9824
rect 17060 9760 17076 9824
rect 17140 9760 17156 9824
rect 17220 9760 17236 9824
rect 17300 9760 17306 9824
rect 16910 9759 17306 9760
rect 22910 9824 23306 9825
rect 22910 9760 22916 9824
rect 22980 9760 22996 9824
rect 23060 9760 23076 9824
rect 23140 9760 23156 9824
rect 23220 9760 23236 9824
rect 23300 9760 23306 9824
rect 22910 9759 23306 9760
rect 28910 9824 29306 9825
rect 28910 9760 28916 9824
rect 28980 9760 28996 9824
rect 29060 9760 29076 9824
rect 29140 9760 29156 9824
rect 29220 9760 29236 9824
rect 29300 9760 29306 9824
rect 28910 9759 29306 9760
rect 4170 9280 4566 9281
rect 4170 9216 4176 9280
rect 4240 9216 4256 9280
rect 4320 9216 4336 9280
rect 4400 9216 4416 9280
rect 4480 9216 4496 9280
rect 4560 9216 4566 9280
rect 4170 9215 4566 9216
rect 10170 9280 10566 9281
rect 10170 9216 10176 9280
rect 10240 9216 10256 9280
rect 10320 9216 10336 9280
rect 10400 9216 10416 9280
rect 10480 9216 10496 9280
rect 10560 9216 10566 9280
rect 10170 9215 10566 9216
rect 16170 9280 16566 9281
rect 16170 9216 16176 9280
rect 16240 9216 16256 9280
rect 16320 9216 16336 9280
rect 16400 9216 16416 9280
rect 16480 9216 16496 9280
rect 16560 9216 16566 9280
rect 16170 9215 16566 9216
rect 22170 9280 22566 9281
rect 22170 9216 22176 9280
rect 22240 9216 22256 9280
rect 22320 9216 22336 9280
rect 22400 9216 22416 9280
rect 22480 9216 22496 9280
rect 22560 9216 22566 9280
rect 22170 9215 22566 9216
rect 28170 9280 28566 9281
rect 28170 9216 28176 9280
rect 28240 9216 28256 9280
rect 28320 9216 28336 9280
rect 28400 9216 28416 9280
rect 28480 9216 28496 9280
rect 28560 9216 28566 9280
rect 28170 9215 28566 9216
rect 10777 8940 10843 8941
rect 10726 8876 10732 8940
rect 10796 8938 10843 8940
rect 10796 8936 10888 8938
rect 10838 8880 10888 8936
rect 10796 8878 10888 8880
rect 10796 8876 10843 8878
rect 10777 8875 10843 8876
rect 4910 8736 5306 8737
rect 4910 8672 4916 8736
rect 4980 8672 4996 8736
rect 5060 8672 5076 8736
rect 5140 8672 5156 8736
rect 5220 8672 5236 8736
rect 5300 8672 5306 8736
rect 4910 8671 5306 8672
rect 10910 8736 11306 8737
rect 10910 8672 10916 8736
rect 10980 8672 10996 8736
rect 11060 8672 11076 8736
rect 11140 8672 11156 8736
rect 11220 8672 11236 8736
rect 11300 8672 11306 8736
rect 10910 8671 11306 8672
rect 16910 8736 17306 8737
rect 16910 8672 16916 8736
rect 16980 8672 16996 8736
rect 17060 8672 17076 8736
rect 17140 8672 17156 8736
rect 17220 8672 17236 8736
rect 17300 8672 17306 8736
rect 16910 8671 17306 8672
rect 22910 8736 23306 8737
rect 22910 8672 22916 8736
rect 22980 8672 22996 8736
rect 23060 8672 23076 8736
rect 23140 8672 23156 8736
rect 23220 8672 23236 8736
rect 23300 8672 23306 8736
rect 22910 8671 23306 8672
rect 28910 8736 29306 8737
rect 28910 8672 28916 8736
rect 28980 8672 28996 8736
rect 29060 8672 29076 8736
rect 29140 8672 29156 8736
rect 29220 8672 29236 8736
rect 29300 8672 29306 8736
rect 28910 8671 29306 8672
rect 10041 8532 10107 8533
rect 9990 8530 9996 8532
rect 9950 8470 9996 8530
rect 10060 8528 10107 8532
rect 10102 8472 10107 8528
rect 9990 8468 9996 8470
rect 10060 8468 10107 8472
rect 10041 8467 10107 8468
rect 14825 8530 14891 8533
rect 26877 8530 26943 8533
rect 14825 8528 26943 8530
rect 14825 8472 14830 8528
rect 14886 8472 26882 8528
rect 26938 8472 26943 8528
rect 14825 8470 26943 8472
rect 14825 8467 14891 8470
rect 26877 8467 26943 8470
rect 4170 8192 4566 8193
rect 4170 8128 4176 8192
rect 4240 8128 4256 8192
rect 4320 8128 4336 8192
rect 4400 8128 4416 8192
rect 4480 8128 4496 8192
rect 4560 8128 4566 8192
rect 4170 8127 4566 8128
rect 10170 8192 10566 8193
rect 10170 8128 10176 8192
rect 10240 8128 10256 8192
rect 10320 8128 10336 8192
rect 10400 8128 10416 8192
rect 10480 8128 10496 8192
rect 10560 8128 10566 8192
rect 10170 8127 10566 8128
rect 16170 8192 16566 8193
rect 16170 8128 16176 8192
rect 16240 8128 16256 8192
rect 16320 8128 16336 8192
rect 16400 8128 16416 8192
rect 16480 8128 16496 8192
rect 16560 8128 16566 8192
rect 16170 8127 16566 8128
rect 22170 8192 22566 8193
rect 22170 8128 22176 8192
rect 22240 8128 22256 8192
rect 22320 8128 22336 8192
rect 22400 8128 22416 8192
rect 22480 8128 22496 8192
rect 22560 8128 22566 8192
rect 22170 8127 22566 8128
rect 28170 8192 28566 8193
rect 28170 8128 28176 8192
rect 28240 8128 28256 8192
rect 28320 8128 28336 8192
rect 28400 8128 28416 8192
rect 28480 8128 28496 8192
rect 28560 8128 28566 8192
rect 28170 8127 28566 8128
rect 4910 7648 5306 7649
rect 4910 7584 4916 7648
rect 4980 7584 4996 7648
rect 5060 7584 5076 7648
rect 5140 7584 5156 7648
rect 5220 7584 5236 7648
rect 5300 7584 5306 7648
rect 4910 7583 5306 7584
rect 10910 7648 11306 7649
rect 10910 7584 10916 7648
rect 10980 7584 10996 7648
rect 11060 7584 11076 7648
rect 11140 7584 11156 7648
rect 11220 7584 11236 7648
rect 11300 7584 11306 7648
rect 10910 7583 11306 7584
rect 16910 7648 17306 7649
rect 16910 7584 16916 7648
rect 16980 7584 16996 7648
rect 17060 7584 17076 7648
rect 17140 7584 17156 7648
rect 17220 7584 17236 7648
rect 17300 7584 17306 7648
rect 16910 7583 17306 7584
rect 22910 7648 23306 7649
rect 22910 7584 22916 7648
rect 22980 7584 22996 7648
rect 23060 7584 23076 7648
rect 23140 7584 23156 7648
rect 23220 7584 23236 7648
rect 23300 7584 23306 7648
rect 22910 7583 23306 7584
rect 28910 7648 29306 7649
rect 28910 7584 28916 7648
rect 28980 7584 28996 7648
rect 29060 7584 29076 7648
rect 29140 7584 29156 7648
rect 29220 7584 29236 7648
rect 29300 7584 29306 7648
rect 28910 7583 29306 7584
rect 31845 7578 31911 7581
rect 32174 7578 32974 7608
rect 31845 7576 32974 7578
rect 31845 7520 31850 7576
rect 31906 7520 32974 7576
rect 31845 7518 32974 7520
rect 31845 7515 31911 7518
rect 32174 7488 32974 7518
rect 9673 7442 9739 7445
rect 9673 7440 9874 7442
rect 9673 7384 9678 7440
rect 9734 7384 9874 7440
rect 9673 7382 9874 7384
rect 9673 7379 9739 7382
rect 9814 7306 9874 7382
rect 15377 7306 15443 7309
rect 9814 7304 15443 7306
rect 9814 7248 15382 7304
rect 15438 7248 15443 7304
rect 9814 7246 15443 7248
rect 15377 7243 15443 7246
rect 4170 7104 4566 7105
rect 4170 7040 4176 7104
rect 4240 7040 4256 7104
rect 4320 7040 4336 7104
rect 4400 7040 4416 7104
rect 4480 7040 4496 7104
rect 4560 7040 4566 7104
rect 4170 7039 4566 7040
rect 10170 7104 10566 7105
rect 10170 7040 10176 7104
rect 10240 7040 10256 7104
rect 10320 7040 10336 7104
rect 10400 7040 10416 7104
rect 10480 7040 10496 7104
rect 10560 7040 10566 7104
rect 10170 7039 10566 7040
rect 16170 7104 16566 7105
rect 16170 7040 16176 7104
rect 16240 7040 16256 7104
rect 16320 7040 16336 7104
rect 16400 7040 16416 7104
rect 16480 7040 16496 7104
rect 16560 7040 16566 7104
rect 16170 7039 16566 7040
rect 22170 7104 22566 7105
rect 22170 7040 22176 7104
rect 22240 7040 22256 7104
rect 22320 7040 22336 7104
rect 22400 7040 22416 7104
rect 22480 7040 22496 7104
rect 22560 7040 22566 7104
rect 22170 7039 22566 7040
rect 28170 7104 28566 7105
rect 28170 7040 28176 7104
rect 28240 7040 28256 7104
rect 28320 7040 28336 7104
rect 28400 7040 28416 7104
rect 28480 7040 28496 7104
rect 28560 7040 28566 7104
rect 28170 7039 28566 7040
rect 9765 6762 9831 6765
rect 10726 6762 10732 6764
rect 9765 6760 10732 6762
rect 9765 6704 9770 6760
rect 9826 6704 10732 6760
rect 9765 6702 10732 6704
rect 9765 6699 9831 6702
rect 10726 6700 10732 6702
rect 10796 6762 10802 6764
rect 17309 6762 17375 6765
rect 10796 6760 17375 6762
rect 10796 6704 17314 6760
rect 17370 6704 17375 6760
rect 10796 6702 17375 6704
rect 10796 6700 10802 6702
rect 17309 6699 17375 6702
rect 4910 6560 5306 6561
rect 4910 6496 4916 6560
rect 4980 6496 4996 6560
rect 5060 6496 5076 6560
rect 5140 6496 5156 6560
rect 5220 6496 5236 6560
rect 5300 6496 5306 6560
rect 4910 6495 5306 6496
rect 10910 6560 11306 6561
rect 10910 6496 10916 6560
rect 10980 6496 10996 6560
rect 11060 6496 11076 6560
rect 11140 6496 11156 6560
rect 11220 6496 11236 6560
rect 11300 6496 11306 6560
rect 10910 6495 11306 6496
rect 16910 6560 17306 6561
rect 16910 6496 16916 6560
rect 16980 6496 16996 6560
rect 17060 6496 17076 6560
rect 17140 6496 17156 6560
rect 17220 6496 17236 6560
rect 17300 6496 17306 6560
rect 16910 6495 17306 6496
rect 22910 6560 23306 6561
rect 22910 6496 22916 6560
rect 22980 6496 22996 6560
rect 23060 6496 23076 6560
rect 23140 6496 23156 6560
rect 23220 6496 23236 6560
rect 23300 6496 23306 6560
rect 22910 6495 23306 6496
rect 28910 6560 29306 6561
rect 28910 6496 28916 6560
rect 28980 6496 28996 6560
rect 29060 6496 29076 6560
rect 29140 6496 29156 6560
rect 29220 6496 29236 6560
rect 29300 6496 29306 6560
rect 28910 6495 29306 6496
rect 0 6218 800 6248
rect 933 6218 999 6221
rect 0 6216 999 6218
rect 0 6160 938 6216
rect 994 6160 999 6216
rect 0 6158 999 6160
rect 0 6128 800 6158
rect 933 6155 999 6158
rect 4170 6016 4566 6017
rect 4170 5952 4176 6016
rect 4240 5952 4256 6016
rect 4320 5952 4336 6016
rect 4400 5952 4416 6016
rect 4480 5952 4496 6016
rect 4560 5952 4566 6016
rect 4170 5951 4566 5952
rect 10170 6016 10566 6017
rect 10170 5952 10176 6016
rect 10240 5952 10256 6016
rect 10320 5952 10336 6016
rect 10400 5952 10416 6016
rect 10480 5952 10496 6016
rect 10560 5952 10566 6016
rect 10170 5951 10566 5952
rect 16170 6016 16566 6017
rect 16170 5952 16176 6016
rect 16240 5952 16256 6016
rect 16320 5952 16336 6016
rect 16400 5952 16416 6016
rect 16480 5952 16496 6016
rect 16560 5952 16566 6016
rect 16170 5951 16566 5952
rect 22170 6016 22566 6017
rect 22170 5952 22176 6016
rect 22240 5952 22256 6016
rect 22320 5952 22336 6016
rect 22400 5952 22416 6016
rect 22480 5952 22496 6016
rect 22560 5952 22566 6016
rect 22170 5951 22566 5952
rect 28170 6016 28566 6017
rect 28170 5952 28176 6016
rect 28240 5952 28256 6016
rect 28320 5952 28336 6016
rect 28400 5952 28416 6016
rect 28480 5952 28496 6016
rect 28560 5952 28566 6016
rect 28170 5951 28566 5952
rect 4910 5472 5306 5473
rect 4910 5408 4916 5472
rect 4980 5408 4996 5472
rect 5060 5408 5076 5472
rect 5140 5408 5156 5472
rect 5220 5408 5236 5472
rect 5300 5408 5306 5472
rect 4910 5407 5306 5408
rect 10910 5472 11306 5473
rect 10910 5408 10916 5472
rect 10980 5408 10996 5472
rect 11060 5408 11076 5472
rect 11140 5408 11156 5472
rect 11220 5408 11236 5472
rect 11300 5408 11306 5472
rect 10910 5407 11306 5408
rect 16910 5472 17306 5473
rect 16910 5408 16916 5472
rect 16980 5408 16996 5472
rect 17060 5408 17076 5472
rect 17140 5408 17156 5472
rect 17220 5408 17236 5472
rect 17300 5408 17306 5472
rect 16910 5407 17306 5408
rect 22910 5472 23306 5473
rect 22910 5408 22916 5472
rect 22980 5408 22996 5472
rect 23060 5408 23076 5472
rect 23140 5408 23156 5472
rect 23220 5408 23236 5472
rect 23300 5408 23306 5472
rect 22910 5407 23306 5408
rect 28910 5472 29306 5473
rect 28910 5408 28916 5472
rect 28980 5408 28996 5472
rect 29060 5408 29076 5472
rect 29140 5408 29156 5472
rect 29220 5408 29236 5472
rect 29300 5408 29306 5472
rect 28910 5407 29306 5408
rect 10041 4996 10107 4997
rect 9990 4994 9996 4996
rect 9950 4934 9996 4994
rect 10060 4992 10107 4996
rect 10102 4936 10107 4992
rect 9990 4932 9996 4934
rect 10060 4932 10107 4936
rect 10041 4931 10107 4932
rect 4170 4928 4566 4929
rect 4170 4864 4176 4928
rect 4240 4864 4256 4928
rect 4320 4864 4336 4928
rect 4400 4864 4416 4928
rect 4480 4864 4496 4928
rect 4560 4864 4566 4928
rect 4170 4863 4566 4864
rect 10170 4928 10566 4929
rect 10170 4864 10176 4928
rect 10240 4864 10256 4928
rect 10320 4864 10336 4928
rect 10400 4864 10416 4928
rect 10480 4864 10496 4928
rect 10560 4864 10566 4928
rect 10170 4863 10566 4864
rect 16170 4928 16566 4929
rect 16170 4864 16176 4928
rect 16240 4864 16256 4928
rect 16320 4864 16336 4928
rect 16400 4864 16416 4928
rect 16480 4864 16496 4928
rect 16560 4864 16566 4928
rect 16170 4863 16566 4864
rect 22170 4928 22566 4929
rect 22170 4864 22176 4928
rect 22240 4864 22256 4928
rect 22320 4864 22336 4928
rect 22400 4864 22416 4928
rect 22480 4864 22496 4928
rect 22560 4864 22566 4928
rect 22170 4863 22566 4864
rect 28170 4928 28566 4929
rect 28170 4864 28176 4928
rect 28240 4864 28256 4928
rect 28320 4864 28336 4928
rect 28400 4864 28416 4928
rect 28480 4864 28496 4928
rect 28560 4864 28566 4928
rect 28170 4863 28566 4864
rect 4910 4384 5306 4385
rect 4910 4320 4916 4384
rect 4980 4320 4996 4384
rect 5060 4320 5076 4384
rect 5140 4320 5156 4384
rect 5220 4320 5236 4384
rect 5300 4320 5306 4384
rect 4910 4319 5306 4320
rect 10910 4384 11306 4385
rect 10910 4320 10916 4384
rect 10980 4320 10996 4384
rect 11060 4320 11076 4384
rect 11140 4320 11156 4384
rect 11220 4320 11236 4384
rect 11300 4320 11306 4384
rect 10910 4319 11306 4320
rect 16910 4384 17306 4385
rect 16910 4320 16916 4384
rect 16980 4320 16996 4384
rect 17060 4320 17076 4384
rect 17140 4320 17156 4384
rect 17220 4320 17236 4384
rect 17300 4320 17306 4384
rect 16910 4319 17306 4320
rect 22910 4384 23306 4385
rect 22910 4320 22916 4384
rect 22980 4320 22996 4384
rect 23060 4320 23076 4384
rect 23140 4320 23156 4384
rect 23220 4320 23236 4384
rect 23300 4320 23306 4384
rect 22910 4319 23306 4320
rect 28910 4384 29306 4385
rect 28910 4320 28916 4384
rect 28980 4320 28996 4384
rect 29060 4320 29076 4384
rect 29140 4320 29156 4384
rect 29220 4320 29236 4384
rect 29300 4320 29306 4384
rect 28910 4319 29306 4320
rect 4170 3840 4566 3841
rect 4170 3776 4176 3840
rect 4240 3776 4256 3840
rect 4320 3776 4336 3840
rect 4400 3776 4416 3840
rect 4480 3776 4496 3840
rect 4560 3776 4566 3840
rect 4170 3775 4566 3776
rect 10170 3840 10566 3841
rect 10170 3776 10176 3840
rect 10240 3776 10256 3840
rect 10320 3776 10336 3840
rect 10400 3776 10416 3840
rect 10480 3776 10496 3840
rect 10560 3776 10566 3840
rect 10170 3775 10566 3776
rect 16170 3840 16566 3841
rect 16170 3776 16176 3840
rect 16240 3776 16256 3840
rect 16320 3776 16336 3840
rect 16400 3776 16416 3840
rect 16480 3776 16496 3840
rect 16560 3776 16566 3840
rect 16170 3775 16566 3776
rect 22170 3840 22566 3841
rect 22170 3776 22176 3840
rect 22240 3776 22256 3840
rect 22320 3776 22336 3840
rect 22400 3776 22416 3840
rect 22480 3776 22496 3840
rect 22560 3776 22566 3840
rect 22170 3775 22566 3776
rect 28170 3840 28566 3841
rect 28170 3776 28176 3840
rect 28240 3776 28256 3840
rect 28320 3776 28336 3840
rect 28400 3776 28416 3840
rect 28480 3776 28496 3840
rect 28560 3776 28566 3840
rect 28170 3775 28566 3776
rect 4910 3296 5306 3297
rect 4910 3232 4916 3296
rect 4980 3232 4996 3296
rect 5060 3232 5076 3296
rect 5140 3232 5156 3296
rect 5220 3232 5236 3296
rect 5300 3232 5306 3296
rect 4910 3231 5306 3232
rect 10910 3296 11306 3297
rect 10910 3232 10916 3296
rect 10980 3232 10996 3296
rect 11060 3232 11076 3296
rect 11140 3232 11156 3296
rect 11220 3232 11236 3296
rect 11300 3232 11306 3296
rect 10910 3231 11306 3232
rect 16910 3296 17306 3297
rect 16910 3232 16916 3296
rect 16980 3232 16996 3296
rect 17060 3232 17076 3296
rect 17140 3232 17156 3296
rect 17220 3232 17236 3296
rect 17300 3232 17306 3296
rect 16910 3231 17306 3232
rect 22910 3296 23306 3297
rect 22910 3232 22916 3296
rect 22980 3232 22996 3296
rect 23060 3232 23076 3296
rect 23140 3232 23156 3296
rect 23220 3232 23236 3296
rect 23300 3232 23306 3296
rect 22910 3231 23306 3232
rect 28910 3296 29306 3297
rect 28910 3232 28916 3296
rect 28980 3232 28996 3296
rect 29060 3232 29076 3296
rect 29140 3232 29156 3296
rect 29220 3232 29236 3296
rect 29300 3232 29306 3296
rect 28910 3231 29306 3232
rect 4170 2752 4566 2753
rect 4170 2688 4176 2752
rect 4240 2688 4256 2752
rect 4320 2688 4336 2752
rect 4400 2688 4416 2752
rect 4480 2688 4496 2752
rect 4560 2688 4566 2752
rect 4170 2687 4566 2688
rect 10170 2752 10566 2753
rect 10170 2688 10176 2752
rect 10240 2688 10256 2752
rect 10320 2688 10336 2752
rect 10400 2688 10416 2752
rect 10480 2688 10496 2752
rect 10560 2688 10566 2752
rect 10170 2687 10566 2688
rect 16170 2752 16566 2753
rect 16170 2688 16176 2752
rect 16240 2688 16256 2752
rect 16320 2688 16336 2752
rect 16400 2688 16416 2752
rect 16480 2688 16496 2752
rect 16560 2688 16566 2752
rect 16170 2687 16566 2688
rect 22170 2752 22566 2753
rect 22170 2688 22176 2752
rect 22240 2688 22256 2752
rect 22320 2688 22336 2752
rect 22400 2688 22416 2752
rect 22480 2688 22496 2752
rect 22560 2688 22566 2752
rect 22170 2687 22566 2688
rect 28170 2752 28566 2753
rect 28170 2688 28176 2752
rect 28240 2688 28256 2752
rect 28320 2688 28336 2752
rect 28400 2688 28416 2752
rect 28480 2688 28496 2752
rect 28560 2688 28566 2752
rect 28170 2687 28566 2688
rect 14038 2484 14044 2548
rect 14108 2546 14114 2548
rect 17033 2546 17099 2549
rect 14108 2544 17099 2546
rect 14108 2488 17038 2544
rect 17094 2488 17099 2544
rect 14108 2486 17099 2488
rect 14108 2484 14114 2486
rect 17033 2483 17099 2486
rect 4910 2208 5306 2209
rect 4910 2144 4916 2208
rect 4980 2144 4996 2208
rect 5060 2144 5076 2208
rect 5140 2144 5156 2208
rect 5220 2144 5236 2208
rect 5300 2144 5306 2208
rect 4910 2143 5306 2144
rect 10910 2208 11306 2209
rect 10910 2144 10916 2208
rect 10980 2144 10996 2208
rect 11060 2144 11076 2208
rect 11140 2144 11156 2208
rect 11220 2144 11236 2208
rect 11300 2144 11306 2208
rect 10910 2143 11306 2144
rect 16910 2208 17306 2209
rect 16910 2144 16916 2208
rect 16980 2144 16996 2208
rect 17060 2144 17076 2208
rect 17140 2144 17156 2208
rect 17220 2144 17236 2208
rect 17300 2144 17306 2208
rect 16910 2143 17306 2144
rect 22910 2208 23306 2209
rect 22910 2144 22916 2208
rect 22980 2144 22996 2208
rect 23060 2144 23076 2208
rect 23140 2144 23156 2208
rect 23220 2144 23236 2208
rect 23300 2144 23306 2208
rect 22910 2143 23306 2144
rect 28910 2208 29306 2209
rect 28910 2144 28916 2208
rect 28980 2144 28996 2208
rect 29060 2144 29076 2208
rect 29140 2144 29156 2208
rect 29220 2144 29236 2208
rect 29300 2144 29306 2208
rect 28910 2143 29306 2144
rect 31385 1458 31451 1461
rect 32174 1458 32974 1488
rect 31385 1456 32974 1458
rect 31385 1400 31390 1456
rect 31446 1400 32974 1456
rect 31385 1398 32974 1400
rect 31385 1395 31451 1398
rect 32174 1368 32974 1398
<< via3 >>
rect 4916 32668 4980 32672
rect 4916 32612 4920 32668
rect 4920 32612 4976 32668
rect 4976 32612 4980 32668
rect 4916 32608 4980 32612
rect 4996 32668 5060 32672
rect 4996 32612 5000 32668
rect 5000 32612 5056 32668
rect 5056 32612 5060 32668
rect 4996 32608 5060 32612
rect 5076 32668 5140 32672
rect 5076 32612 5080 32668
rect 5080 32612 5136 32668
rect 5136 32612 5140 32668
rect 5076 32608 5140 32612
rect 5156 32668 5220 32672
rect 5156 32612 5160 32668
rect 5160 32612 5216 32668
rect 5216 32612 5220 32668
rect 5156 32608 5220 32612
rect 5236 32668 5300 32672
rect 5236 32612 5240 32668
rect 5240 32612 5296 32668
rect 5296 32612 5300 32668
rect 5236 32608 5300 32612
rect 10916 32668 10980 32672
rect 10916 32612 10920 32668
rect 10920 32612 10976 32668
rect 10976 32612 10980 32668
rect 10916 32608 10980 32612
rect 10996 32668 11060 32672
rect 10996 32612 11000 32668
rect 11000 32612 11056 32668
rect 11056 32612 11060 32668
rect 10996 32608 11060 32612
rect 11076 32668 11140 32672
rect 11076 32612 11080 32668
rect 11080 32612 11136 32668
rect 11136 32612 11140 32668
rect 11076 32608 11140 32612
rect 11156 32668 11220 32672
rect 11156 32612 11160 32668
rect 11160 32612 11216 32668
rect 11216 32612 11220 32668
rect 11156 32608 11220 32612
rect 11236 32668 11300 32672
rect 11236 32612 11240 32668
rect 11240 32612 11296 32668
rect 11296 32612 11300 32668
rect 11236 32608 11300 32612
rect 16916 32668 16980 32672
rect 16916 32612 16920 32668
rect 16920 32612 16976 32668
rect 16976 32612 16980 32668
rect 16916 32608 16980 32612
rect 16996 32668 17060 32672
rect 16996 32612 17000 32668
rect 17000 32612 17056 32668
rect 17056 32612 17060 32668
rect 16996 32608 17060 32612
rect 17076 32668 17140 32672
rect 17076 32612 17080 32668
rect 17080 32612 17136 32668
rect 17136 32612 17140 32668
rect 17076 32608 17140 32612
rect 17156 32668 17220 32672
rect 17156 32612 17160 32668
rect 17160 32612 17216 32668
rect 17216 32612 17220 32668
rect 17156 32608 17220 32612
rect 17236 32668 17300 32672
rect 17236 32612 17240 32668
rect 17240 32612 17296 32668
rect 17296 32612 17300 32668
rect 17236 32608 17300 32612
rect 22916 32668 22980 32672
rect 22916 32612 22920 32668
rect 22920 32612 22976 32668
rect 22976 32612 22980 32668
rect 22916 32608 22980 32612
rect 22996 32668 23060 32672
rect 22996 32612 23000 32668
rect 23000 32612 23056 32668
rect 23056 32612 23060 32668
rect 22996 32608 23060 32612
rect 23076 32668 23140 32672
rect 23076 32612 23080 32668
rect 23080 32612 23136 32668
rect 23136 32612 23140 32668
rect 23076 32608 23140 32612
rect 23156 32668 23220 32672
rect 23156 32612 23160 32668
rect 23160 32612 23216 32668
rect 23216 32612 23220 32668
rect 23156 32608 23220 32612
rect 23236 32668 23300 32672
rect 23236 32612 23240 32668
rect 23240 32612 23296 32668
rect 23296 32612 23300 32668
rect 23236 32608 23300 32612
rect 28916 32668 28980 32672
rect 28916 32612 28920 32668
rect 28920 32612 28976 32668
rect 28976 32612 28980 32668
rect 28916 32608 28980 32612
rect 28996 32668 29060 32672
rect 28996 32612 29000 32668
rect 29000 32612 29056 32668
rect 29056 32612 29060 32668
rect 28996 32608 29060 32612
rect 29076 32668 29140 32672
rect 29076 32612 29080 32668
rect 29080 32612 29136 32668
rect 29136 32612 29140 32668
rect 29076 32608 29140 32612
rect 29156 32668 29220 32672
rect 29156 32612 29160 32668
rect 29160 32612 29216 32668
rect 29216 32612 29220 32668
rect 29156 32608 29220 32612
rect 29236 32668 29300 32672
rect 29236 32612 29240 32668
rect 29240 32612 29296 32668
rect 29296 32612 29300 32668
rect 29236 32608 29300 32612
rect 4176 32124 4240 32128
rect 4176 32068 4180 32124
rect 4180 32068 4236 32124
rect 4236 32068 4240 32124
rect 4176 32064 4240 32068
rect 4256 32124 4320 32128
rect 4256 32068 4260 32124
rect 4260 32068 4316 32124
rect 4316 32068 4320 32124
rect 4256 32064 4320 32068
rect 4336 32124 4400 32128
rect 4336 32068 4340 32124
rect 4340 32068 4396 32124
rect 4396 32068 4400 32124
rect 4336 32064 4400 32068
rect 4416 32124 4480 32128
rect 4416 32068 4420 32124
rect 4420 32068 4476 32124
rect 4476 32068 4480 32124
rect 4416 32064 4480 32068
rect 4496 32124 4560 32128
rect 4496 32068 4500 32124
rect 4500 32068 4556 32124
rect 4556 32068 4560 32124
rect 4496 32064 4560 32068
rect 10176 32124 10240 32128
rect 10176 32068 10180 32124
rect 10180 32068 10236 32124
rect 10236 32068 10240 32124
rect 10176 32064 10240 32068
rect 10256 32124 10320 32128
rect 10256 32068 10260 32124
rect 10260 32068 10316 32124
rect 10316 32068 10320 32124
rect 10256 32064 10320 32068
rect 10336 32124 10400 32128
rect 10336 32068 10340 32124
rect 10340 32068 10396 32124
rect 10396 32068 10400 32124
rect 10336 32064 10400 32068
rect 10416 32124 10480 32128
rect 10416 32068 10420 32124
rect 10420 32068 10476 32124
rect 10476 32068 10480 32124
rect 10416 32064 10480 32068
rect 10496 32124 10560 32128
rect 10496 32068 10500 32124
rect 10500 32068 10556 32124
rect 10556 32068 10560 32124
rect 10496 32064 10560 32068
rect 16176 32124 16240 32128
rect 16176 32068 16180 32124
rect 16180 32068 16236 32124
rect 16236 32068 16240 32124
rect 16176 32064 16240 32068
rect 16256 32124 16320 32128
rect 16256 32068 16260 32124
rect 16260 32068 16316 32124
rect 16316 32068 16320 32124
rect 16256 32064 16320 32068
rect 16336 32124 16400 32128
rect 16336 32068 16340 32124
rect 16340 32068 16396 32124
rect 16396 32068 16400 32124
rect 16336 32064 16400 32068
rect 16416 32124 16480 32128
rect 16416 32068 16420 32124
rect 16420 32068 16476 32124
rect 16476 32068 16480 32124
rect 16416 32064 16480 32068
rect 16496 32124 16560 32128
rect 16496 32068 16500 32124
rect 16500 32068 16556 32124
rect 16556 32068 16560 32124
rect 16496 32064 16560 32068
rect 22176 32124 22240 32128
rect 22176 32068 22180 32124
rect 22180 32068 22236 32124
rect 22236 32068 22240 32124
rect 22176 32064 22240 32068
rect 22256 32124 22320 32128
rect 22256 32068 22260 32124
rect 22260 32068 22316 32124
rect 22316 32068 22320 32124
rect 22256 32064 22320 32068
rect 22336 32124 22400 32128
rect 22336 32068 22340 32124
rect 22340 32068 22396 32124
rect 22396 32068 22400 32124
rect 22336 32064 22400 32068
rect 22416 32124 22480 32128
rect 22416 32068 22420 32124
rect 22420 32068 22476 32124
rect 22476 32068 22480 32124
rect 22416 32064 22480 32068
rect 22496 32124 22560 32128
rect 22496 32068 22500 32124
rect 22500 32068 22556 32124
rect 22556 32068 22560 32124
rect 22496 32064 22560 32068
rect 28176 32124 28240 32128
rect 28176 32068 28180 32124
rect 28180 32068 28236 32124
rect 28236 32068 28240 32124
rect 28176 32064 28240 32068
rect 28256 32124 28320 32128
rect 28256 32068 28260 32124
rect 28260 32068 28316 32124
rect 28316 32068 28320 32124
rect 28256 32064 28320 32068
rect 28336 32124 28400 32128
rect 28336 32068 28340 32124
rect 28340 32068 28396 32124
rect 28396 32068 28400 32124
rect 28336 32064 28400 32068
rect 28416 32124 28480 32128
rect 28416 32068 28420 32124
rect 28420 32068 28476 32124
rect 28476 32068 28480 32124
rect 28416 32064 28480 32068
rect 28496 32124 28560 32128
rect 28496 32068 28500 32124
rect 28500 32068 28556 32124
rect 28556 32068 28560 32124
rect 28496 32064 28560 32068
rect 27844 31860 27908 31924
rect 4916 31580 4980 31584
rect 4916 31524 4920 31580
rect 4920 31524 4976 31580
rect 4976 31524 4980 31580
rect 4916 31520 4980 31524
rect 4996 31580 5060 31584
rect 4996 31524 5000 31580
rect 5000 31524 5056 31580
rect 5056 31524 5060 31580
rect 4996 31520 5060 31524
rect 5076 31580 5140 31584
rect 5076 31524 5080 31580
rect 5080 31524 5136 31580
rect 5136 31524 5140 31580
rect 5076 31520 5140 31524
rect 5156 31580 5220 31584
rect 5156 31524 5160 31580
rect 5160 31524 5216 31580
rect 5216 31524 5220 31580
rect 5156 31520 5220 31524
rect 5236 31580 5300 31584
rect 5236 31524 5240 31580
rect 5240 31524 5296 31580
rect 5296 31524 5300 31580
rect 5236 31520 5300 31524
rect 10916 31580 10980 31584
rect 10916 31524 10920 31580
rect 10920 31524 10976 31580
rect 10976 31524 10980 31580
rect 10916 31520 10980 31524
rect 10996 31580 11060 31584
rect 10996 31524 11000 31580
rect 11000 31524 11056 31580
rect 11056 31524 11060 31580
rect 10996 31520 11060 31524
rect 11076 31580 11140 31584
rect 11076 31524 11080 31580
rect 11080 31524 11136 31580
rect 11136 31524 11140 31580
rect 11076 31520 11140 31524
rect 11156 31580 11220 31584
rect 11156 31524 11160 31580
rect 11160 31524 11216 31580
rect 11216 31524 11220 31580
rect 11156 31520 11220 31524
rect 11236 31580 11300 31584
rect 11236 31524 11240 31580
rect 11240 31524 11296 31580
rect 11296 31524 11300 31580
rect 11236 31520 11300 31524
rect 16916 31580 16980 31584
rect 16916 31524 16920 31580
rect 16920 31524 16976 31580
rect 16976 31524 16980 31580
rect 16916 31520 16980 31524
rect 16996 31580 17060 31584
rect 16996 31524 17000 31580
rect 17000 31524 17056 31580
rect 17056 31524 17060 31580
rect 16996 31520 17060 31524
rect 17076 31580 17140 31584
rect 17076 31524 17080 31580
rect 17080 31524 17136 31580
rect 17136 31524 17140 31580
rect 17076 31520 17140 31524
rect 17156 31580 17220 31584
rect 17156 31524 17160 31580
rect 17160 31524 17216 31580
rect 17216 31524 17220 31580
rect 17156 31520 17220 31524
rect 17236 31580 17300 31584
rect 17236 31524 17240 31580
rect 17240 31524 17296 31580
rect 17296 31524 17300 31580
rect 17236 31520 17300 31524
rect 22916 31580 22980 31584
rect 22916 31524 22920 31580
rect 22920 31524 22976 31580
rect 22976 31524 22980 31580
rect 22916 31520 22980 31524
rect 22996 31580 23060 31584
rect 22996 31524 23000 31580
rect 23000 31524 23056 31580
rect 23056 31524 23060 31580
rect 22996 31520 23060 31524
rect 23076 31580 23140 31584
rect 23076 31524 23080 31580
rect 23080 31524 23136 31580
rect 23136 31524 23140 31580
rect 23076 31520 23140 31524
rect 23156 31580 23220 31584
rect 23156 31524 23160 31580
rect 23160 31524 23216 31580
rect 23216 31524 23220 31580
rect 23156 31520 23220 31524
rect 23236 31580 23300 31584
rect 23236 31524 23240 31580
rect 23240 31524 23296 31580
rect 23296 31524 23300 31580
rect 23236 31520 23300 31524
rect 28916 31580 28980 31584
rect 28916 31524 28920 31580
rect 28920 31524 28976 31580
rect 28976 31524 28980 31580
rect 28916 31520 28980 31524
rect 28996 31580 29060 31584
rect 28996 31524 29000 31580
rect 29000 31524 29056 31580
rect 29056 31524 29060 31580
rect 28996 31520 29060 31524
rect 29076 31580 29140 31584
rect 29076 31524 29080 31580
rect 29080 31524 29136 31580
rect 29136 31524 29140 31580
rect 29076 31520 29140 31524
rect 29156 31580 29220 31584
rect 29156 31524 29160 31580
rect 29160 31524 29216 31580
rect 29216 31524 29220 31580
rect 29156 31520 29220 31524
rect 29236 31580 29300 31584
rect 29236 31524 29240 31580
rect 29240 31524 29296 31580
rect 29296 31524 29300 31580
rect 29236 31520 29300 31524
rect 4176 31036 4240 31040
rect 4176 30980 4180 31036
rect 4180 30980 4236 31036
rect 4236 30980 4240 31036
rect 4176 30976 4240 30980
rect 4256 31036 4320 31040
rect 4256 30980 4260 31036
rect 4260 30980 4316 31036
rect 4316 30980 4320 31036
rect 4256 30976 4320 30980
rect 4336 31036 4400 31040
rect 4336 30980 4340 31036
rect 4340 30980 4396 31036
rect 4396 30980 4400 31036
rect 4336 30976 4400 30980
rect 4416 31036 4480 31040
rect 4416 30980 4420 31036
rect 4420 30980 4476 31036
rect 4476 30980 4480 31036
rect 4416 30976 4480 30980
rect 4496 31036 4560 31040
rect 4496 30980 4500 31036
rect 4500 30980 4556 31036
rect 4556 30980 4560 31036
rect 4496 30976 4560 30980
rect 10176 31036 10240 31040
rect 10176 30980 10180 31036
rect 10180 30980 10236 31036
rect 10236 30980 10240 31036
rect 10176 30976 10240 30980
rect 10256 31036 10320 31040
rect 10256 30980 10260 31036
rect 10260 30980 10316 31036
rect 10316 30980 10320 31036
rect 10256 30976 10320 30980
rect 10336 31036 10400 31040
rect 10336 30980 10340 31036
rect 10340 30980 10396 31036
rect 10396 30980 10400 31036
rect 10336 30976 10400 30980
rect 10416 31036 10480 31040
rect 10416 30980 10420 31036
rect 10420 30980 10476 31036
rect 10476 30980 10480 31036
rect 10416 30976 10480 30980
rect 10496 31036 10560 31040
rect 10496 30980 10500 31036
rect 10500 30980 10556 31036
rect 10556 30980 10560 31036
rect 10496 30976 10560 30980
rect 16176 31036 16240 31040
rect 16176 30980 16180 31036
rect 16180 30980 16236 31036
rect 16236 30980 16240 31036
rect 16176 30976 16240 30980
rect 16256 31036 16320 31040
rect 16256 30980 16260 31036
rect 16260 30980 16316 31036
rect 16316 30980 16320 31036
rect 16256 30976 16320 30980
rect 16336 31036 16400 31040
rect 16336 30980 16340 31036
rect 16340 30980 16396 31036
rect 16396 30980 16400 31036
rect 16336 30976 16400 30980
rect 16416 31036 16480 31040
rect 16416 30980 16420 31036
rect 16420 30980 16476 31036
rect 16476 30980 16480 31036
rect 16416 30976 16480 30980
rect 16496 31036 16560 31040
rect 16496 30980 16500 31036
rect 16500 30980 16556 31036
rect 16556 30980 16560 31036
rect 16496 30976 16560 30980
rect 22176 31036 22240 31040
rect 22176 30980 22180 31036
rect 22180 30980 22236 31036
rect 22236 30980 22240 31036
rect 22176 30976 22240 30980
rect 22256 31036 22320 31040
rect 22256 30980 22260 31036
rect 22260 30980 22316 31036
rect 22316 30980 22320 31036
rect 22256 30976 22320 30980
rect 22336 31036 22400 31040
rect 22336 30980 22340 31036
rect 22340 30980 22396 31036
rect 22396 30980 22400 31036
rect 22336 30976 22400 30980
rect 22416 31036 22480 31040
rect 22416 30980 22420 31036
rect 22420 30980 22476 31036
rect 22476 30980 22480 31036
rect 22416 30976 22480 30980
rect 22496 31036 22560 31040
rect 22496 30980 22500 31036
rect 22500 30980 22556 31036
rect 22556 30980 22560 31036
rect 22496 30976 22560 30980
rect 28176 31036 28240 31040
rect 28176 30980 28180 31036
rect 28180 30980 28236 31036
rect 28236 30980 28240 31036
rect 28176 30976 28240 30980
rect 28256 31036 28320 31040
rect 28256 30980 28260 31036
rect 28260 30980 28316 31036
rect 28316 30980 28320 31036
rect 28256 30976 28320 30980
rect 28336 31036 28400 31040
rect 28336 30980 28340 31036
rect 28340 30980 28396 31036
rect 28396 30980 28400 31036
rect 28336 30976 28400 30980
rect 28416 31036 28480 31040
rect 28416 30980 28420 31036
rect 28420 30980 28476 31036
rect 28476 30980 28480 31036
rect 28416 30976 28480 30980
rect 28496 31036 28560 31040
rect 28496 30980 28500 31036
rect 28500 30980 28556 31036
rect 28556 30980 28560 31036
rect 28496 30976 28560 30980
rect 4916 30492 4980 30496
rect 4916 30436 4920 30492
rect 4920 30436 4976 30492
rect 4976 30436 4980 30492
rect 4916 30432 4980 30436
rect 4996 30492 5060 30496
rect 4996 30436 5000 30492
rect 5000 30436 5056 30492
rect 5056 30436 5060 30492
rect 4996 30432 5060 30436
rect 5076 30492 5140 30496
rect 5076 30436 5080 30492
rect 5080 30436 5136 30492
rect 5136 30436 5140 30492
rect 5076 30432 5140 30436
rect 5156 30492 5220 30496
rect 5156 30436 5160 30492
rect 5160 30436 5216 30492
rect 5216 30436 5220 30492
rect 5156 30432 5220 30436
rect 5236 30492 5300 30496
rect 5236 30436 5240 30492
rect 5240 30436 5296 30492
rect 5296 30436 5300 30492
rect 5236 30432 5300 30436
rect 10916 30492 10980 30496
rect 10916 30436 10920 30492
rect 10920 30436 10976 30492
rect 10976 30436 10980 30492
rect 10916 30432 10980 30436
rect 10996 30492 11060 30496
rect 10996 30436 11000 30492
rect 11000 30436 11056 30492
rect 11056 30436 11060 30492
rect 10996 30432 11060 30436
rect 11076 30492 11140 30496
rect 11076 30436 11080 30492
rect 11080 30436 11136 30492
rect 11136 30436 11140 30492
rect 11076 30432 11140 30436
rect 11156 30492 11220 30496
rect 11156 30436 11160 30492
rect 11160 30436 11216 30492
rect 11216 30436 11220 30492
rect 11156 30432 11220 30436
rect 11236 30492 11300 30496
rect 11236 30436 11240 30492
rect 11240 30436 11296 30492
rect 11296 30436 11300 30492
rect 11236 30432 11300 30436
rect 16916 30492 16980 30496
rect 16916 30436 16920 30492
rect 16920 30436 16976 30492
rect 16976 30436 16980 30492
rect 16916 30432 16980 30436
rect 16996 30492 17060 30496
rect 16996 30436 17000 30492
rect 17000 30436 17056 30492
rect 17056 30436 17060 30492
rect 16996 30432 17060 30436
rect 17076 30492 17140 30496
rect 17076 30436 17080 30492
rect 17080 30436 17136 30492
rect 17136 30436 17140 30492
rect 17076 30432 17140 30436
rect 17156 30492 17220 30496
rect 17156 30436 17160 30492
rect 17160 30436 17216 30492
rect 17216 30436 17220 30492
rect 17156 30432 17220 30436
rect 17236 30492 17300 30496
rect 17236 30436 17240 30492
rect 17240 30436 17296 30492
rect 17296 30436 17300 30492
rect 17236 30432 17300 30436
rect 22916 30492 22980 30496
rect 22916 30436 22920 30492
rect 22920 30436 22976 30492
rect 22976 30436 22980 30492
rect 22916 30432 22980 30436
rect 22996 30492 23060 30496
rect 22996 30436 23000 30492
rect 23000 30436 23056 30492
rect 23056 30436 23060 30492
rect 22996 30432 23060 30436
rect 23076 30492 23140 30496
rect 23076 30436 23080 30492
rect 23080 30436 23136 30492
rect 23136 30436 23140 30492
rect 23076 30432 23140 30436
rect 23156 30492 23220 30496
rect 23156 30436 23160 30492
rect 23160 30436 23216 30492
rect 23216 30436 23220 30492
rect 23156 30432 23220 30436
rect 23236 30492 23300 30496
rect 23236 30436 23240 30492
rect 23240 30436 23296 30492
rect 23296 30436 23300 30492
rect 23236 30432 23300 30436
rect 28916 30492 28980 30496
rect 28916 30436 28920 30492
rect 28920 30436 28976 30492
rect 28976 30436 28980 30492
rect 28916 30432 28980 30436
rect 28996 30492 29060 30496
rect 28996 30436 29000 30492
rect 29000 30436 29056 30492
rect 29056 30436 29060 30492
rect 28996 30432 29060 30436
rect 29076 30492 29140 30496
rect 29076 30436 29080 30492
rect 29080 30436 29136 30492
rect 29136 30436 29140 30492
rect 29076 30432 29140 30436
rect 29156 30492 29220 30496
rect 29156 30436 29160 30492
rect 29160 30436 29216 30492
rect 29216 30436 29220 30492
rect 29156 30432 29220 30436
rect 29236 30492 29300 30496
rect 29236 30436 29240 30492
rect 29240 30436 29296 30492
rect 29296 30436 29300 30492
rect 29236 30432 29300 30436
rect 4176 29948 4240 29952
rect 4176 29892 4180 29948
rect 4180 29892 4236 29948
rect 4236 29892 4240 29948
rect 4176 29888 4240 29892
rect 4256 29948 4320 29952
rect 4256 29892 4260 29948
rect 4260 29892 4316 29948
rect 4316 29892 4320 29948
rect 4256 29888 4320 29892
rect 4336 29948 4400 29952
rect 4336 29892 4340 29948
rect 4340 29892 4396 29948
rect 4396 29892 4400 29948
rect 4336 29888 4400 29892
rect 4416 29948 4480 29952
rect 4416 29892 4420 29948
rect 4420 29892 4476 29948
rect 4476 29892 4480 29948
rect 4416 29888 4480 29892
rect 4496 29948 4560 29952
rect 4496 29892 4500 29948
rect 4500 29892 4556 29948
rect 4556 29892 4560 29948
rect 4496 29888 4560 29892
rect 10176 29948 10240 29952
rect 10176 29892 10180 29948
rect 10180 29892 10236 29948
rect 10236 29892 10240 29948
rect 10176 29888 10240 29892
rect 10256 29948 10320 29952
rect 10256 29892 10260 29948
rect 10260 29892 10316 29948
rect 10316 29892 10320 29948
rect 10256 29888 10320 29892
rect 10336 29948 10400 29952
rect 10336 29892 10340 29948
rect 10340 29892 10396 29948
rect 10396 29892 10400 29948
rect 10336 29888 10400 29892
rect 10416 29948 10480 29952
rect 10416 29892 10420 29948
rect 10420 29892 10476 29948
rect 10476 29892 10480 29948
rect 10416 29888 10480 29892
rect 10496 29948 10560 29952
rect 10496 29892 10500 29948
rect 10500 29892 10556 29948
rect 10556 29892 10560 29948
rect 10496 29888 10560 29892
rect 16176 29948 16240 29952
rect 16176 29892 16180 29948
rect 16180 29892 16236 29948
rect 16236 29892 16240 29948
rect 16176 29888 16240 29892
rect 16256 29948 16320 29952
rect 16256 29892 16260 29948
rect 16260 29892 16316 29948
rect 16316 29892 16320 29948
rect 16256 29888 16320 29892
rect 16336 29948 16400 29952
rect 16336 29892 16340 29948
rect 16340 29892 16396 29948
rect 16396 29892 16400 29948
rect 16336 29888 16400 29892
rect 16416 29948 16480 29952
rect 16416 29892 16420 29948
rect 16420 29892 16476 29948
rect 16476 29892 16480 29948
rect 16416 29888 16480 29892
rect 16496 29948 16560 29952
rect 16496 29892 16500 29948
rect 16500 29892 16556 29948
rect 16556 29892 16560 29948
rect 16496 29888 16560 29892
rect 22176 29948 22240 29952
rect 22176 29892 22180 29948
rect 22180 29892 22236 29948
rect 22236 29892 22240 29948
rect 22176 29888 22240 29892
rect 22256 29948 22320 29952
rect 22256 29892 22260 29948
rect 22260 29892 22316 29948
rect 22316 29892 22320 29948
rect 22256 29888 22320 29892
rect 22336 29948 22400 29952
rect 22336 29892 22340 29948
rect 22340 29892 22396 29948
rect 22396 29892 22400 29948
rect 22336 29888 22400 29892
rect 22416 29948 22480 29952
rect 22416 29892 22420 29948
rect 22420 29892 22476 29948
rect 22476 29892 22480 29948
rect 22416 29888 22480 29892
rect 22496 29948 22560 29952
rect 22496 29892 22500 29948
rect 22500 29892 22556 29948
rect 22556 29892 22560 29948
rect 22496 29888 22560 29892
rect 28176 29948 28240 29952
rect 28176 29892 28180 29948
rect 28180 29892 28236 29948
rect 28236 29892 28240 29948
rect 28176 29888 28240 29892
rect 28256 29948 28320 29952
rect 28256 29892 28260 29948
rect 28260 29892 28316 29948
rect 28316 29892 28320 29948
rect 28256 29888 28320 29892
rect 28336 29948 28400 29952
rect 28336 29892 28340 29948
rect 28340 29892 28396 29948
rect 28396 29892 28400 29948
rect 28336 29888 28400 29892
rect 28416 29948 28480 29952
rect 28416 29892 28420 29948
rect 28420 29892 28476 29948
rect 28476 29892 28480 29948
rect 28416 29888 28480 29892
rect 28496 29948 28560 29952
rect 28496 29892 28500 29948
rect 28500 29892 28556 29948
rect 28556 29892 28560 29948
rect 28496 29888 28560 29892
rect 4916 29404 4980 29408
rect 4916 29348 4920 29404
rect 4920 29348 4976 29404
rect 4976 29348 4980 29404
rect 4916 29344 4980 29348
rect 4996 29404 5060 29408
rect 4996 29348 5000 29404
rect 5000 29348 5056 29404
rect 5056 29348 5060 29404
rect 4996 29344 5060 29348
rect 5076 29404 5140 29408
rect 5076 29348 5080 29404
rect 5080 29348 5136 29404
rect 5136 29348 5140 29404
rect 5076 29344 5140 29348
rect 5156 29404 5220 29408
rect 5156 29348 5160 29404
rect 5160 29348 5216 29404
rect 5216 29348 5220 29404
rect 5156 29344 5220 29348
rect 5236 29404 5300 29408
rect 5236 29348 5240 29404
rect 5240 29348 5296 29404
rect 5296 29348 5300 29404
rect 5236 29344 5300 29348
rect 10916 29404 10980 29408
rect 10916 29348 10920 29404
rect 10920 29348 10976 29404
rect 10976 29348 10980 29404
rect 10916 29344 10980 29348
rect 10996 29404 11060 29408
rect 10996 29348 11000 29404
rect 11000 29348 11056 29404
rect 11056 29348 11060 29404
rect 10996 29344 11060 29348
rect 11076 29404 11140 29408
rect 11076 29348 11080 29404
rect 11080 29348 11136 29404
rect 11136 29348 11140 29404
rect 11076 29344 11140 29348
rect 11156 29404 11220 29408
rect 11156 29348 11160 29404
rect 11160 29348 11216 29404
rect 11216 29348 11220 29404
rect 11156 29344 11220 29348
rect 11236 29404 11300 29408
rect 11236 29348 11240 29404
rect 11240 29348 11296 29404
rect 11296 29348 11300 29404
rect 11236 29344 11300 29348
rect 16916 29404 16980 29408
rect 16916 29348 16920 29404
rect 16920 29348 16976 29404
rect 16976 29348 16980 29404
rect 16916 29344 16980 29348
rect 16996 29404 17060 29408
rect 16996 29348 17000 29404
rect 17000 29348 17056 29404
rect 17056 29348 17060 29404
rect 16996 29344 17060 29348
rect 17076 29404 17140 29408
rect 17076 29348 17080 29404
rect 17080 29348 17136 29404
rect 17136 29348 17140 29404
rect 17076 29344 17140 29348
rect 17156 29404 17220 29408
rect 17156 29348 17160 29404
rect 17160 29348 17216 29404
rect 17216 29348 17220 29404
rect 17156 29344 17220 29348
rect 17236 29404 17300 29408
rect 17236 29348 17240 29404
rect 17240 29348 17296 29404
rect 17296 29348 17300 29404
rect 17236 29344 17300 29348
rect 22916 29404 22980 29408
rect 22916 29348 22920 29404
rect 22920 29348 22976 29404
rect 22976 29348 22980 29404
rect 22916 29344 22980 29348
rect 22996 29404 23060 29408
rect 22996 29348 23000 29404
rect 23000 29348 23056 29404
rect 23056 29348 23060 29404
rect 22996 29344 23060 29348
rect 23076 29404 23140 29408
rect 23076 29348 23080 29404
rect 23080 29348 23136 29404
rect 23136 29348 23140 29404
rect 23076 29344 23140 29348
rect 23156 29404 23220 29408
rect 23156 29348 23160 29404
rect 23160 29348 23216 29404
rect 23216 29348 23220 29404
rect 23156 29344 23220 29348
rect 23236 29404 23300 29408
rect 23236 29348 23240 29404
rect 23240 29348 23296 29404
rect 23296 29348 23300 29404
rect 23236 29344 23300 29348
rect 28916 29404 28980 29408
rect 28916 29348 28920 29404
rect 28920 29348 28976 29404
rect 28976 29348 28980 29404
rect 28916 29344 28980 29348
rect 28996 29404 29060 29408
rect 28996 29348 29000 29404
rect 29000 29348 29056 29404
rect 29056 29348 29060 29404
rect 28996 29344 29060 29348
rect 29076 29404 29140 29408
rect 29076 29348 29080 29404
rect 29080 29348 29136 29404
rect 29136 29348 29140 29404
rect 29076 29344 29140 29348
rect 29156 29404 29220 29408
rect 29156 29348 29160 29404
rect 29160 29348 29216 29404
rect 29216 29348 29220 29404
rect 29156 29344 29220 29348
rect 29236 29404 29300 29408
rect 29236 29348 29240 29404
rect 29240 29348 29296 29404
rect 29296 29348 29300 29404
rect 29236 29344 29300 29348
rect 14044 29064 14108 29068
rect 14044 29008 14058 29064
rect 14058 29008 14108 29064
rect 14044 29004 14108 29008
rect 4176 28860 4240 28864
rect 4176 28804 4180 28860
rect 4180 28804 4236 28860
rect 4236 28804 4240 28860
rect 4176 28800 4240 28804
rect 4256 28860 4320 28864
rect 4256 28804 4260 28860
rect 4260 28804 4316 28860
rect 4316 28804 4320 28860
rect 4256 28800 4320 28804
rect 4336 28860 4400 28864
rect 4336 28804 4340 28860
rect 4340 28804 4396 28860
rect 4396 28804 4400 28860
rect 4336 28800 4400 28804
rect 4416 28860 4480 28864
rect 4416 28804 4420 28860
rect 4420 28804 4476 28860
rect 4476 28804 4480 28860
rect 4416 28800 4480 28804
rect 4496 28860 4560 28864
rect 4496 28804 4500 28860
rect 4500 28804 4556 28860
rect 4556 28804 4560 28860
rect 4496 28800 4560 28804
rect 10176 28860 10240 28864
rect 10176 28804 10180 28860
rect 10180 28804 10236 28860
rect 10236 28804 10240 28860
rect 10176 28800 10240 28804
rect 10256 28860 10320 28864
rect 10256 28804 10260 28860
rect 10260 28804 10316 28860
rect 10316 28804 10320 28860
rect 10256 28800 10320 28804
rect 10336 28860 10400 28864
rect 10336 28804 10340 28860
rect 10340 28804 10396 28860
rect 10396 28804 10400 28860
rect 10336 28800 10400 28804
rect 10416 28860 10480 28864
rect 10416 28804 10420 28860
rect 10420 28804 10476 28860
rect 10476 28804 10480 28860
rect 10416 28800 10480 28804
rect 10496 28860 10560 28864
rect 10496 28804 10500 28860
rect 10500 28804 10556 28860
rect 10556 28804 10560 28860
rect 10496 28800 10560 28804
rect 16176 28860 16240 28864
rect 16176 28804 16180 28860
rect 16180 28804 16236 28860
rect 16236 28804 16240 28860
rect 16176 28800 16240 28804
rect 16256 28860 16320 28864
rect 16256 28804 16260 28860
rect 16260 28804 16316 28860
rect 16316 28804 16320 28860
rect 16256 28800 16320 28804
rect 16336 28860 16400 28864
rect 16336 28804 16340 28860
rect 16340 28804 16396 28860
rect 16396 28804 16400 28860
rect 16336 28800 16400 28804
rect 16416 28860 16480 28864
rect 16416 28804 16420 28860
rect 16420 28804 16476 28860
rect 16476 28804 16480 28860
rect 16416 28800 16480 28804
rect 16496 28860 16560 28864
rect 16496 28804 16500 28860
rect 16500 28804 16556 28860
rect 16556 28804 16560 28860
rect 16496 28800 16560 28804
rect 22176 28860 22240 28864
rect 22176 28804 22180 28860
rect 22180 28804 22236 28860
rect 22236 28804 22240 28860
rect 22176 28800 22240 28804
rect 22256 28860 22320 28864
rect 22256 28804 22260 28860
rect 22260 28804 22316 28860
rect 22316 28804 22320 28860
rect 22256 28800 22320 28804
rect 22336 28860 22400 28864
rect 22336 28804 22340 28860
rect 22340 28804 22396 28860
rect 22396 28804 22400 28860
rect 22336 28800 22400 28804
rect 22416 28860 22480 28864
rect 22416 28804 22420 28860
rect 22420 28804 22476 28860
rect 22476 28804 22480 28860
rect 22416 28800 22480 28804
rect 22496 28860 22560 28864
rect 22496 28804 22500 28860
rect 22500 28804 22556 28860
rect 22556 28804 22560 28860
rect 22496 28800 22560 28804
rect 28176 28860 28240 28864
rect 28176 28804 28180 28860
rect 28180 28804 28236 28860
rect 28236 28804 28240 28860
rect 28176 28800 28240 28804
rect 28256 28860 28320 28864
rect 28256 28804 28260 28860
rect 28260 28804 28316 28860
rect 28316 28804 28320 28860
rect 28256 28800 28320 28804
rect 28336 28860 28400 28864
rect 28336 28804 28340 28860
rect 28340 28804 28396 28860
rect 28396 28804 28400 28860
rect 28336 28800 28400 28804
rect 28416 28860 28480 28864
rect 28416 28804 28420 28860
rect 28420 28804 28476 28860
rect 28476 28804 28480 28860
rect 28416 28800 28480 28804
rect 28496 28860 28560 28864
rect 28496 28804 28500 28860
rect 28500 28804 28556 28860
rect 28556 28804 28560 28860
rect 28496 28800 28560 28804
rect 4916 28316 4980 28320
rect 4916 28260 4920 28316
rect 4920 28260 4976 28316
rect 4976 28260 4980 28316
rect 4916 28256 4980 28260
rect 4996 28316 5060 28320
rect 4996 28260 5000 28316
rect 5000 28260 5056 28316
rect 5056 28260 5060 28316
rect 4996 28256 5060 28260
rect 5076 28316 5140 28320
rect 5076 28260 5080 28316
rect 5080 28260 5136 28316
rect 5136 28260 5140 28316
rect 5076 28256 5140 28260
rect 5156 28316 5220 28320
rect 5156 28260 5160 28316
rect 5160 28260 5216 28316
rect 5216 28260 5220 28316
rect 5156 28256 5220 28260
rect 5236 28316 5300 28320
rect 5236 28260 5240 28316
rect 5240 28260 5296 28316
rect 5296 28260 5300 28316
rect 5236 28256 5300 28260
rect 10916 28316 10980 28320
rect 10916 28260 10920 28316
rect 10920 28260 10976 28316
rect 10976 28260 10980 28316
rect 10916 28256 10980 28260
rect 10996 28316 11060 28320
rect 10996 28260 11000 28316
rect 11000 28260 11056 28316
rect 11056 28260 11060 28316
rect 10996 28256 11060 28260
rect 11076 28316 11140 28320
rect 11076 28260 11080 28316
rect 11080 28260 11136 28316
rect 11136 28260 11140 28316
rect 11076 28256 11140 28260
rect 11156 28316 11220 28320
rect 11156 28260 11160 28316
rect 11160 28260 11216 28316
rect 11216 28260 11220 28316
rect 11156 28256 11220 28260
rect 11236 28316 11300 28320
rect 11236 28260 11240 28316
rect 11240 28260 11296 28316
rect 11296 28260 11300 28316
rect 11236 28256 11300 28260
rect 16916 28316 16980 28320
rect 16916 28260 16920 28316
rect 16920 28260 16976 28316
rect 16976 28260 16980 28316
rect 16916 28256 16980 28260
rect 16996 28316 17060 28320
rect 16996 28260 17000 28316
rect 17000 28260 17056 28316
rect 17056 28260 17060 28316
rect 16996 28256 17060 28260
rect 17076 28316 17140 28320
rect 17076 28260 17080 28316
rect 17080 28260 17136 28316
rect 17136 28260 17140 28316
rect 17076 28256 17140 28260
rect 17156 28316 17220 28320
rect 17156 28260 17160 28316
rect 17160 28260 17216 28316
rect 17216 28260 17220 28316
rect 17156 28256 17220 28260
rect 17236 28316 17300 28320
rect 17236 28260 17240 28316
rect 17240 28260 17296 28316
rect 17296 28260 17300 28316
rect 17236 28256 17300 28260
rect 22916 28316 22980 28320
rect 22916 28260 22920 28316
rect 22920 28260 22976 28316
rect 22976 28260 22980 28316
rect 22916 28256 22980 28260
rect 22996 28316 23060 28320
rect 22996 28260 23000 28316
rect 23000 28260 23056 28316
rect 23056 28260 23060 28316
rect 22996 28256 23060 28260
rect 23076 28316 23140 28320
rect 23076 28260 23080 28316
rect 23080 28260 23136 28316
rect 23136 28260 23140 28316
rect 23076 28256 23140 28260
rect 23156 28316 23220 28320
rect 23156 28260 23160 28316
rect 23160 28260 23216 28316
rect 23216 28260 23220 28316
rect 23156 28256 23220 28260
rect 23236 28316 23300 28320
rect 23236 28260 23240 28316
rect 23240 28260 23296 28316
rect 23296 28260 23300 28316
rect 23236 28256 23300 28260
rect 28916 28316 28980 28320
rect 28916 28260 28920 28316
rect 28920 28260 28976 28316
rect 28976 28260 28980 28316
rect 28916 28256 28980 28260
rect 28996 28316 29060 28320
rect 28996 28260 29000 28316
rect 29000 28260 29056 28316
rect 29056 28260 29060 28316
rect 28996 28256 29060 28260
rect 29076 28316 29140 28320
rect 29076 28260 29080 28316
rect 29080 28260 29136 28316
rect 29136 28260 29140 28316
rect 29076 28256 29140 28260
rect 29156 28316 29220 28320
rect 29156 28260 29160 28316
rect 29160 28260 29216 28316
rect 29216 28260 29220 28316
rect 29156 28256 29220 28260
rect 29236 28316 29300 28320
rect 29236 28260 29240 28316
rect 29240 28260 29296 28316
rect 29296 28260 29300 28316
rect 29236 28256 29300 28260
rect 4176 27772 4240 27776
rect 4176 27716 4180 27772
rect 4180 27716 4236 27772
rect 4236 27716 4240 27772
rect 4176 27712 4240 27716
rect 4256 27772 4320 27776
rect 4256 27716 4260 27772
rect 4260 27716 4316 27772
rect 4316 27716 4320 27772
rect 4256 27712 4320 27716
rect 4336 27772 4400 27776
rect 4336 27716 4340 27772
rect 4340 27716 4396 27772
rect 4396 27716 4400 27772
rect 4336 27712 4400 27716
rect 4416 27772 4480 27776
rect 4416 27716 4420 27772
rect 4420 27716 4476 27772
rect 4476 27716 4480 27772
rect 4416 27712 4480 27716
rect 4496 27772 4560 27776
rect 4496 27716 4500 27772
rect 4500 27716 4556 27772
rect 4556 27716 4560 27772
rect 4496 27712 4560 27716
rect 10176 27772 10240 27776
rect 10176 27716 10180 27772
rect 10180 27716 10236 27772
rect 10236 27716 10240 27772
rect 10176 27712 10240 27716
rect 10256 27772 10320 27776
rect 10256 27716 10260 27772
rect 10260 27716 10316 27772
rect 10316 27716 10320 27772
rect 10256 27712 10320 27716
rect 10336 27772 10400 27776
rect 10336 27716 10340 27772
rect 10340 27716 10396 27772
rect 10396 27716 10400 27772
rect 10336 27712 10400 27716
rect 10416 27772 10480 27776
rect 10416 27716 10420 27772
rect 10420 27716 10476 27772
rect 10476 27716 10480 27772
rect 10416 27712 10480 27716
rect 10496 27772 10560 27776
rect 10496 27716 10500 27772
rect 10500 27716 10556 27772
rect 10556 27716 10560 27772
rect 10496 27712 10560 27716
rect 16176 27772 16240 27776
rect 16176 27716 16180 27772
rect 16180 27716 16236 27772
rect 16236 27716 16240 27772
rect 16176 27712 16240 27716
rect 16256 27772 16320 27776
rect 16256 27716 16260 27772
rect 16260 27716 16316 27772
rect 16316 27716 16320 27772
rect 16256 27712 16320 27716
rect 16336 27772 16400 27776
rect 16336 27716 16340 27772
rect 16340 27716 16396 27772
rect 16396 27716 16400 27772
rect 16336 27712 16400 27716
rect 16416 27772 16480 27776
rect 16416 27716 16420 27772
rect 16420 27716 16476 27772
rect 16476 27716 16480 27772
rect 16416 27712 16480 27716
rect 16496 27772 16560 27776
rect 16496 27716 16500 27772
rect 16500 27716 16556 27772
rect 16556 27716 16560 27772
rect 16496 27712 16560 27716
rect 22176 27772 22240 27776
rect 22176 27716 22180 27772
rect 22180 27716 22236 27772
rect 22236 27716 22240 27772
rect 22176 27712 22240 27716
rect 22256 27772 22320 27776
rect 22256 27716 22260 27772
rect 22260 27716 22316 27772
rect 22316 27716 22320 27772
rect 22256 27712 22320 27716
rect 22336 27772 22400 27776
rect 22336 27716 22340 27772
rect 22340 27716 22396 27772
rect 22396 27716 22400 27772
rect 22336 27712 22400 27716
rect 22416 27772 22480 27776
rect 22416 27716 22420 27772
rect 22420 27716 22476 27772
rect 22476 27716 22480 27772
rect 22416 27712 22480 27716
rect 22496 27772 22560 27776
rect 22496 27716 22500 27772
rect 22500 27716 22556 27772
rect 22556 27716 22560 27772
rect 22496 27712 22560 27716
rect 28176 27772 28240 27776
rect 28176 27716 28180 27772
rect 28180 27716 28236 27772
rect 28236 27716 28240 27772
rect 28176 27712 28240 27716
rect 28256 27772 28320 27776
rect 28256 27716 28260 27772
rect 28260 27716 28316 27772
rect 28316 27716 28320 27772
rect 28256 27712 28320 27716
rect 28336 27772 28400 27776
rect 28336 27716 28340 27772
rect 28340 27716 28396 27772
rect 28396 27716 28400 27772
rect 28336 27712 28400 27716
rect 28416 27772 28480 27776
rect 28416 27716 28420 27772
rect 28420 27716 28476 27772
rect 28476 27716 28480 27772
rect 28416 27712 28480 27716
rect 28496 27772 28560 27776
rect 28496 27716 28500 27772
rect 28500 27716 28556 27772
rect 28556 27716 28560 27772
rect 28496 27712 28560 27716
rect 4916 27228 4980 27232
rect 4916 27172 4920 27228
rect 4920 27172 4976 27228
rect 4976 27172 4980 27228
rect 4916 27168 4980 27172
rect 4996 27228 5060 27232
rect 4996 27172 5000 27228
rect 5000 27172 5056 27228
rect 5056 27172 5060 27228
rect 4996 27168 5060 27172
rect 5076 27228 5140 27232
rect 5076 27172 5080 27228
rect 5080 27172 5136 27228
rect 5136 27172 5140 27228
rect 5076 27168 5140 27172
rect 5156 27228 5220 27232
rect 5156 27172 5160 27228
rect 5160 27172 5216 27228
rect 5216 27172 5220 27228
rect 5156 27168 5220 27172
rect 5236 27228 5300 27232
rect 5236 27172 5240 27228
rect 5240 27172 5296 27228
rect 5296 27172 5300 27228
rect 5236 27168 5300 27172
rect 10916 27228 10980 27232
rect 10916 27172 10920 27228
rect 10920 27172 10976 27228
rect 10976 27172 10980 27228
rect 10916 27168 10980 27172
rect 10996 27228 11060 27232
rect 10996 27172 11000 27228
rect 11000 27172 11056 27228
rect 11056 27172 11060 27228
rect 10996 27168 11060 27172
rect 11076 27228 11140 27232
rect 11076 27172 11080 27228
rect 11080 27172 11136 27228
rect 11136 27172 11140 27228
rect 11076 27168 11140 27172
rect 11156 27228 11220 27232
rect 11156 27172 11160 27228
rect 11160 27172 11216 27228
rect 11216 27172 11220 27228
rect 11156 27168 11220 27172
rect 11236 27228 11300 27232
rect 11236 27172 11240 27228
rect 11240 27172 11296 27228
rect 11296 27172 11300 27228
rect 11236 27168 11300 27172
rect 16916 27228 16980 27232
rect 16916 27172 16920 27228
rect 16920 27172 16976 27228
rect 16976 27172 16980 27228
rect 16916 27168 16980 27172
rect 16996 27228 17060 27232
rect 16996 27172 17000 27228
rect 17000 27172 17056 27228
rect 17056 27172 17060 27228
rect 16996 27168 17060 27172
rect 17076 27228 17140 27232
rect 17076 27172 17080 27228
rect 17080 27172 17136 27228
rect 17136 27172 17140 27228
rect 17076 27168 17140 27172
rect 17156 27228 17220 27232
rect 17156 27172 17160 27228
rect 17160 27172 17216 27228
rect 17216 27172 17220 27228
rect 17156 27168 17220 27172
rect 17236 27228 17300 27232
rect 17236 27172 17240 27228
rect 17240 27172 17296 27228
rect 17296 27172 17300 27228
rect 17236 27168 17300 27172
rect 22916 27228 22980 27232
rect 22916 27172 22920 27228
rect 22920 27172 22976 27228
rect 22976 27172 22980 27228
rect 22916 27168 22980 27172
rect 22996 27228 23060 27232
rect 22996 27172 23000 27228
rect 23000 27172 23056 27228
rect 23056 27172 23060 27228
rect 22996 27168 23060 27172
rect 23076 27228 23140 27232
rect 23076 27172 23080 27228
rect 23080 27172 23136 27228
rect 23136 27172 23140 27228
rect 23076 27168 23140 27172
rect 23156 27228 23220 27232
rect 23156 27172 23160 27228
rect 23160 27172 23216 27228
rect 23216 27172 23220 27228
rect 23156 27168 23220 27172
rect 23236 27228 23300 27232
rect 23236 27172 23240 27228
rect 23240 27172 23296 27228
rect 23296 27172 23300 27228
rect 23236 27168 23300 27172
rect 28916 27228 28980 27232
rect 28916 27172 28920 27228
rect 28920 27172 28976 27228
rect 28976 27172 28980 27228
rect 28916 27168 28980 27172
rect 28996 27228 29060 27232
rect 28996 27172 29000 27228
rect 29000 27172 29056 27228
rect 29056 27172 29060 27228
rect 28996 27168 29060 27172
rect 29076 27228 29140 27232
rect 29076 27172 29080 27228
rect 29080 27172 29136 27228
rect 29136 27172 29140 27228
rect 29076 27168 29140 27172
rect 29156 27228 29220 27232
rect 29156 27172 29160 27228
rect 29160 27172 29216 27228
rect 29216 27172 29220 27228
rect 29156 27168 29220 27172
rect 29236 27228 29300 27232
rect 29236 27172 29240 27228
rect 29240 27172 29296 27228
rect 29296 27172 29300 27228
rect 29236 27168 29300 27172
rect 4176 26684 4240 26688
rect 4176 26628 4180 26684
rect 4180 26628 4236 26684
rect 4236 26628 4240 26684
rect 4176 26624 4240 26628
rect 4256 26684 4320 26688
rect 4256 26628 4260 26684
rect 4260 26628 4316 26684
rect 4316 26628 4320 26684
rect 4256 26624 4320 26628
rect 4336 26684 4400 26688
rect 4336 26628 4340 26684
rect 4340 26628 4396 26684
rect 4396 26628 4400 26684
rect 4336 26624 4400 26628
rect 4416 26684 4480 26688
rect 4416 26628 4420 26684
rect 4420 26628 4476 26684
rect 4476 26628 4480 26684
rect 4416 26624 4480 26628
rect 4496 26684 4560 26688
rect 4496 26628 4500 26684
rect 4500 26628 4556 26684
rect 4556 26628 4560 26684
rect 4496 26624 4560 26628
rect 10176 26684 10240 26688
rect 10176 26628 10180 26684
rect 10180 26628 10236 26684
rect 10236 26628 10240 26684
rect 10176 26624 10240 26628
rect 10256 26684 10320 26688
rect 10256 26628 10260 26684
rect 10260 26628 10316 26684
rect 10316 26628 10320 26684
rect 10256 26624 10320 26628
rect 10336 26684 10400 26688
rect 10336 26628 10340 26684
rect 10340 26628 10396 26684
rect 10396 26628 10400 26684
rect 10336 26624 10400 26628
rect 10416 26684 10480 26688
rect 10416 26628 10420 26684
rect 10420 26628 10476 26684
rect 10476 26628 10480 26684
rect 10416 26624 10480 26628
rect 10496 26684 10560 26688
rect 10496 26628 10500 26684
rect 10500 26628 10556 26684
rect 10556 26628 10560 26684
rect 10496 26624 10560 26628
rect 16176 26684 16240 26688
rect 16176 26628 16180 26684
rect 16180 26628 16236 26684
rect 16236 26628 16240 26684
rect 16176 26624 16240 26628
rect 16256 26684 16320 26688
rect 16256 26628 16260 26684
rect 16260 26628 16316 26684
rect 16316 26628 16320 26684
rect 16256 26624 16320 26628
rect 16336 26684 16400 26688
rect 16336 26628 16340 26684
rect 16340 26628 16396 26684
rect 16396 26628 16400 26684
rect 16336 26624 16400 26628
rect 16416 26684 16480 26688
rect 16416 26628 16420 26684
rect 16420 26628 16476 26684
rect 16476 26628 16480 26684
rect 16416 26624 16480 26628
rect 16496 26684 16560 26688
rect 16496 26628 16500 26684
rect 16500 26628 16556 26684
rect 16556 26628 16560 26684
rect 16496 26624 16560 26628
rect 22176 26684 22240 26688
rect 22176 26628 22180 26684
rect 22180 26628 22236 26684
rect 22236 26628 22240 26684
rect 22176 26624 22240 26628
rect 22256 26684 22320 26688
rect 22256 26628 22260 26684
rect 22260 26628 22316 26684
rect 22316 26628 22320 26684
rect 22256 26624 22320 26628
rect 22336 26684 22400 26688
rect 22336 26628 22340 26684
rect 22340 26628 22396 26684
rect 22396 26628 22400 26684
rect 22336 26624 22400 26628
rect 22416 26684 22480 26688
rect 22416 26628 22420 26684
rect 22420 26628 22476 26684
rect 22476 26628 22480 26684
rect 22416 26624 22480 26628
rect 22496 26684 22560 26688
rect 22496 26628 22500 26684
rect 22500 26628 22556 26684
rect 22556 26628 22560 26684
rect 22496 26624 22560 26628
rect 28176 26684 28240 26688
rect 28176 26628 28180 26684
rect 28180 26628 28236 26684
rect 28236 26628 28240 26684
rect 28176 26624 28240 26628
rect 28256 26684 28320 26688
rect 28256 26628 28260 26684
rect 28260 26628 28316 26684
rect 28316 26628 28320 26684
rect 28256 26624 28320 26628
rect 28336 26684 28400 26688
rect 28336 26628 28340 26684
rect 28340 26628 28396 26684
rect 28396 26628 28400 26684
rect 28336 26624 28400 26628
rect 28416 26684 28480 26688
rect 28416 26628 28420 26684
rect 28420 26628 28476 26684
rect 28476 26628 28480 26684
rect 28416 26624 28480 26628
rect 28496 26684 28560 26688
rect 28496 26628 28500 26684
rect 28500 26628 28556 26684
rect 28556 26628 28560 26684
rect 28496 26624 28560 26628
rect 4916 26140 4980 26144
rect 4916 26084 4920 26140
rect 4920 26084 4976 26140
rect 4976 26084 4980 26140
rect 4916 26080 4980 26084
rect 4996 26140 5060 26144
rect 4996 26084 5000 26140
rect 5000 26084 5056 26140
rect 5056 26084 5060 26140
rect 4996 26080 5060 26084
rect 5076 26140 5140 26144
rect 5076 26084 5080 26140
rect 5080 26084 5136 26140
rect 5136 26084 5140 26140
rect 5076 26080 5140 26084
rect 5156 26140 5220 26144
rect 5156 26084 5160 26140
rect 5160 26084 5216 26140
rect 5216 26084 5220 26140
rect 5156 26080 5220 26084
rect 5236 26140 5300 26144
rect 5236 26084 5240 26140
rect 5240 26084 5296 26140
rect 5296 26084 5300 26140
rect 5236 26080 5300 26084
rect 10916 26140 10980 26144
rect 10916 26084 10920 26140
rect 10920 26084 10976 26140
rect 10976 26084 10980 26140
rect 10916 26080 10980 26084
rect 10996 26140 11060 26144
rect 10996 26084 11000 26140
rect 11000 26084 11056 26140
rect 11056 26084 11060 26140
rect 10996 26080 11060 26084
rect 11076 26140 11140 26144
rect 11076 26084 11080 26140
rect 11080 26084 11136 26140
rect 11136 26084 11140 26140
rect 11076 26080 11140 26084
rect 11156 26140 11220 26144
rect 11156 26084 11160 26140
rect 11160 26084 11216 26140
rect 11216 26084 11220 26140
rect 11156 26080 11220 26084
rect 11236 26140 11300 26144
rect 11236 26084 11240 26140
rect 11240 26084 11296 26140
rect 11296 26084 11300 26140
rect 11236 26080 11300 26084
rect 16916 26140 16980 26144
rect 16916 26084 16920 26140
rect 16920 26084 16976 26140
rect 16976 26084 16980 26140
rect 16916 26080 16980 26084
rect 16996 26140 17060 26144
rect 16996 26084 17000 26140
rect 17000 26084 17056 26140
rect 17056 26084 17060 26140
rect 16996 26080 17060 26084
rect 17076 26140 17140 26144
rect 17076 26084 17080 26140
rect 17080 26084 17136 26140
rect 17136 26084 17140 26140
rect 17076 26080 17140 26084
rect 17156 26140 17220 26144
rect 17156 26084 17160 26140
rect 17160 26084 17216 26140
rect 17216 26084 17220 26140
rect 17156 26080 17220 26084
rect 17236 26140 17300 26144
rect 17236 26084 17240 26140
rect 17240 26084 17296 26140
rect 17296 26084 17300 26140
rect 17236 26080 17300 26084
rect 22916 26140 22980 26144
rect 22916 26084 22920 26140
rect 22920 26084 22976 26140
rect 22976 26084 22980 26140
rect 22916 26080 22980 26084
rect 22996 26140 23060 26144
rect 22996 26084 23000 26140
rect 23000 26084 23056 26140
rect 23056 26084 23060 26140
rect 22996 26080 23060 26084
rect 23076 26140 23140 26144
rect 23076 26084 23080 26140
rect 23080 26084 23136 26140
rect 23136 26084 23140 26140
rect 23076 26080 23140 26084
rect 23156 26140 23220 26144
rect 23156 26084 23160 26140
rect 23160 26084 23216 26140
rect 23216 26084 23220 26140
rect 23156 26080 23220 26084
rect 23236 26140 23300 26144
rect 23236 26084 23240 26140
rect 23240 26084 23296 26140
rect 23296 26084 23300 26140
rect 23236 26080 23300 26084
rect 28916 26140 28980 26144
rect 28916 26084 28920 26140
rect 28920 26084 28976 26140
rect 28976 26084 28980 26140
rect 28916 26080 28980 26084
rect 28996 26140 29060 26144
rect 28996 26084 29000 26140
rect 29000 26084 29056 26140
rect 29056 26084 29060 26140
rect 28996 26080 29060 26084
rect 29076 26140 29140 26144
rect 29076 26084 29080 26140
rect 29080 26084 29136 26140
rect 29136 26084 29140 26140
rect 29076 26080 29140 26084
rect 29156 26140 29220 26144
rect 29156 26084 29160 26140
rect 29160 26084 29216 26140
rect 29216 26084 29220 26140
rect 29156 26080 29220 26084
rect 29236 26140 29300 26144
rect 29236 26084 29240 26140
rect 29240 26084 29296 26140
rect 29296 26084 29300 26140
rect 29236 26080 29300 26084
rect 4176 25596 4240 25600
rect 4176 25540 4180 25596
rect 4180 25540 4236 25596
rect 4236 25540 4240 25596
rect 4176 25536 4240 25540
rect 4256 25596 4320 25600
rect 4256 25540 4260 25596
rect 4260 25540 4316 25596
rect 4316 25540 4320 25596
rect 4256 25536 4320 25540
rect 4336 25596 4400 25600
rect 4336 25540 4340 25596
rect 4340 25540 4396 25596
rect 4396 25540 4400 25596
rect 4336 25536 4400 25540
rect 4416 25596 4480 25600
rect 4416 25540 4420 25596
rect 4420 25540 4476 25596
rect 4476 25540 4480 25596
rect 4416 25536 4480 25540
rect 4496 25596 4560 25600
rect 4496 25540 4500 25596
rect 4500 25540 4556 25596
rect 4556 25540 4560 25596
rect 4496 25536 4560 25540
rect 10176 25596 10240 25600
rect 10176 25540 10180 25596
rect 10180 25540 10236 25596
rect 10236 25540 10240 25596
rect 10176 25536 10240 25540
rect 10256 25596 10320 25600
rect 10256 25540 10260 25596
rect 10260 25540 10316 25596
rect 10316 25540 10320 25596
rect 10256 25536 10320 25540
rect 10336 25596 10400 25600
rect 10336 25540 10340 25596
rect 10340 25540 10396 25596
rect 10396 25540 10400 25596
rect 10336 25536 10400 25540
rect 10416 25596 10480 25600
rect 10416 25540 10420 25596
rect 10420 25540 10476 25596
rect 10476 25540 10480 25596
rect 10416 25536 10480 25540
rect 10496 25596 10560 25600
rect 10496 25540 10500 25596
rect 10500 25540 10556 25596
rect 10556 25540 10560 25596
rect 10496 25536 10560 25540
rect 16176 25596 16240 25600
rect 16176 25540 16180 25596
rect 16180 25540 16236 25596
rect 16236 25540 16240 25596
rect 16176 25536 16240 25540
rect 16256 25596 16320 25600
rect 16256 25540 16260 25596
rect 16260 25540 16316 25596
rect 16316 25540 16320 25596
rect 16256 25536 16320 25540
rect 16336 25596 16400 25600
rect 16336 25540 16340 25596
rect 16340 25540 16396 25596
rect 16396 25540 16400 25596
rect 16336 25536 16400 25540
rect 16416 25596 16480 25600
rect 16416 25540 16420 25596
rect 16420 25540 16476 25596
rect 16476 25540 16480 25596
rect 16416 25536 16480 25540
rect 16496 25596 16560 25600
rect 16496 25540 16500 25596
rect 16500 25540 16556 25596
rect 16556 25540 16560 25596
rect 16496 25536 16560 25540
rect 22176 25596 22240 25600
rect 22176 25540 22180 25596
rect 22180 25540 22236 25596
rect 22236 25540 22240 25596
rect 22176 25536 22240 25540
rect 22256 25596 22320 25600
rect 22256 25540 22260 25596
rect 22260 25540 22316 25596
rect 22316 25540 22320 25596
rect 22256 25536 22320 25540
rect 22336 25596 22400 25600
rect 22336 25540 22340 25596
rect 22340 25540 22396 25596
rect 22396 25540 22400 25596
rect 22336 25536 22400 25540
rect 22416 25596 22480 25600
rect 22416 25540 22420 25596
rect 22420 25540 22476 25596
rect 22476 25540 22480 25596
rect 22416 25536 22480 25540
rect 22496 25596 22560 25600
rect 22496 25540 22500 25596
rect 22500 25540 22556 25596
rect 22556 25540 22560 25596
rect 22496 25536 22560 25540
rect 28176 25596 28240 25600
rect 28176 25540 28180 25596
rect 28180 25540 28236 25596
rect 28236 25540 28240 25596
rect 28176 25536 28240 25540
rect 28256 25596 28320 25600
rect 28256 25540 28260 25596
rect 28260 25540 28316 25596
rect 28316 25540 28320 25596
rect 28256 25536 28320 25540
rect 28336 25596 28400 25600
rect 28336 25540 28340 25596
rect 28340 25540 28396 25596
rect 28396 25540 28400 25596
rect 28336 25536 28400 25540
rect 28416 25596 28480 25600
rect 28416 25540 28420 25596
rect 28420 25540 28476 25596
rect 28476 25540 28480 25596
rect 28416 25536 28480 25540
rect 28496 25596 28560 25600
rect 28496 25540 28500 25596
rect 28500 25540 28556 25596
rect 28556 25540 28560 25596
rect 28496 25536 28560 25540
rect 4916 25052 4980 25056
rect 4916 24996 4920 25052
rect 4920 24996 4976 25052
rect 4976 24996 4980 25052
rect 4916 24992 4980 24996
rect 4996 25052 5060 25056
rect 4996 24996 5000 25052
rect 5000 24996 5056 25052
rect 5056 24996 5060 25052
rect 4996 24992 5060 24996
rect 5076 25052 5140 25056
rect 5076 24996 5080 25052
rect 5080 24996 5136 25052
rect 5136 24996 5140 25052
rect 5076 24992 5140 24996
rect 5156 25052 5220 25056
rect 5156 24996 5160 25052
rect 5160 24996 5216 25052
rect 5216 24996 5220 25052
rect 5156 24992 5220 24996
rect 5236 25052 5300 25056
rect 5236 24996 5240 25052
rect 5240 24996 5296 25052
rect 5296 24996 5300 25052
rect 5236 24992 5300 24996
rect 10916 25052 10980 25056
rect 10916 24996 10920 25052
rect 10920 24996 10976 25052
rect 10976 24996 10980 25052
rect 10916 24992 10980 24996
rect 10996 25052 11060 25056
rect 10996 24996 11000 25052
rect 11000 24996 11056 25052
rect 11056 24996 11060 25052
rect 10996 24992 11060 24996
rect 11076 25052 11140 25056
rect 11076 24996 11080 25052
rect 11080 24996 11136 25052
rect 11136 24996 11140 25052
rect 11076 24992 11140 24996
rect 11156 25052 11220 25056
rect 11156 24996 11160 25052
rect 11160 24996 11216 25052
rect 11216 24996 11220 25052
rect 11156 24992 11220 24996
rect 11236 25052 11300 25056
rect 11236 24996 11240 25052
rect 11240 24996 11296 25052
rect 11296 24996 11300 25052
rect 11236 24992 11300 24996
rect 16916 25052 16980 25056
rect 16916 24996 16920 25052
rect 16920 24996 16976 25052
rect 16976 24996 16980 25052
rect 16916 24992 16980 24996
rect 16996 25052 17060 25056
rect 16996 24996 17000 25052
rect 17000 24996 17056 25052
rect 17056 24996 17060 25052
rect 16996 24992 17060 24996
rect 17076 25052 17140 25056
rect 17076 24996 17080 25052
rect 17080 24996 17136 25052
rect 17136 24996 17140 25052
rect 17076 24992 17140 24996
rect 17156 25052 17220 25056
rect 17156 24996 17160 25052
rect 17160 24996 17216 25052
rect 17216 24996 17220 25052
rect 17156 24992 17220 24996
rect 17236 25052 17300 25056
rect 17236 24996 17240 25052
rect 17240 24996 17296 25052
rect 17296 24996 17300 25052
rect 17236 24992 17300 24996
rect 22916 25052 22980 25056
rect 22916 24996 22920 25052
rect 22920 24996 22976 25052
rect 22976 24996 22980 25052
rect 22916 24992 22980 24996
rect 22996 25052 23060 25056
rect 22996 24996 23000 25052
rect 23000 24996 23056 25052
rect 23056 24996 23060 25052
rect 22996 24992 23060 24996
rect 23076 25052 23140 25056
rect 23076 24996 23080 25052
rect 23080 24996 23136 25052
rect 23136 24996 23140 25052
rect 23076 24992 23140 24996
rect 23156 25052 23220 25056
rect 23156 24996 23160 25052
rect 23160 24996 23216 25052
rect 23216 24996 23220 25052
rect 23156 24992 23220 24996
rect 23236 25052 23300 25056
rect 23236 24996 23240 25052
rect 23240 24996 23296 25052
rect 23296 24996 23300 25052
rect 23236 24992 23300 24996
rect 28916 25052 28980 25056
rect 28916 24996 28920 25052
rect 28920 24996 28976 25052
rect 28976 24996 28980 25052
rect 28916 24992 28980 24996
rect 28996 25052 29060 25056
rect 28996 24996 29000 25052
rect 29000 24996 29056 25052
rect 29056 24996 29060 25052
rect 28996 24992 29060 24996
rect 29076 25052 29140 25056
rect 29076 24996 29080 25052
rect 29080 24996 29136 25052
rect 29136 24996 29140 25052
rect 29076 24992 29140 24996
rect 29156 25052 29220 25056
rect 29156 24996 29160 25052
rect 29160 24996 29216 25052
rect 29216 24996 29220 25052
rect 29156 24992 29220 24996
rect 29236 25052 29300 25056
rect 29236 24996 29240 25052
rect 29240 24996 29296 25052
rect 29296 24996 29300 25052
rect 29236 24992 29300 24996
rect 4176 24508 4240 24512
rect 4176 24452 4180 24508
rect 4180 24452 4236 24508
rect 4236 24452 4240 24508
rect 4176 24448 4240 24452
rect 4256 24508 4320 24512
rect 4256 24452 4260 24508
rect 4260 24452 4316 24508
rect 4316 24452 4320 24508
rect 4256 24448 4320 24452
rect 4336 24508 4400 24512
rect 4336 24452 4340 24508
rect 4340 24452 4396 24508
rect 4396 24452 4400 24508
rect 4336 24448 4400 24452
rect 4416 24508 4480 24512
rect 4416 24452 4420 24508
rect 4420 24452 4476 24508
rect 4476 24452 4480 24508
rect 4416 24448 4480 24452
rect 4496 24508 4560 24512
rect 4496 24452 4500 24508
rect 4500 24452 4556 24508
rect 4556 24452 4560 24508
rect 4496 24448 4560 24452
rect 10176 24508 10240 24512
rect 10176 24452 10180 24508
rect 10180 24452 10236 24508
rect 10236 24452 10240 24508
rect 10176 24448 10240 24452
rect 10256 24508 10320 24512
rect 10256 24452 10260 24508
rect 10260 24452 10316 24508
rect 10316 24452 10320 24508
rect 10256 24448 10320 24452
rect 10336 24508 10400 24512
rect 10336 24452 10340 24508
rect 10340 24452 10396 24508
rect 10396 24452 10400 24508
rect 10336 24448 10400 24452
rect 10416 24508 10480 24512
rect 10416 24452 10420 24508
rect 10420 24452 10476 24508
rect 10476 24452 10480 24508
rect 10416 24448 10480 24452
rect 10496 24508 10560 24512
rect 10496 24452 10500 24508
rect 10500 24452 10556 24508
rect 10556 24452 10560 24508
rect 10496 24448 10560 24452
rect 16176 24508 16240 24512
rect 16176 24452 16180 24508
rect 16180 24452 16236 24508
rect 16236 24452 16240 24508
rect 16176 24448 16240 24452
rect 16256 24508 16320 24512
rect 16256 24452 16260 24508
rect 16260 24452 16316 24508
rect 16316 24452 16320 24508
rect 16256 24448 16320 24452
rect 16336 24508 16400 24512
rect 16336 24452 16340 24508
rect 16340 24452 16396 24508
rect 16396 24452 16400 24508
rect 16336 24448 16400 24452
rect 16416 24508 16480 24512
rect 16416 24452 16420 24508
rect 16420 24452 16476 24508
rect 16476 24452 16480 24508
rect 16416 24448 16480 24452
rect 16496 24508 16560 24512
rect 16496 24452 16500 24508
rect 16500 24452 16556 24508
rect 16556 24452 16560 24508
rect 16496 24448 16560 24452
rect 22176 24508 22240 24512
rect 22176 24452 22180 24508
rect 22180 24452 22236 24508
rect 22236 24452 22240 24508
rect 22176 24448 22240 24452
rect 22256 24508 22320 24512
rect 22256 24452 22260 24508
rect 22260 24452 22316 24508
rect 22316 24452 22320 24508
rect 22256 24448 22320 24452
rect 22336 24508 22400 24512
rect 22336 24452 22340 24508
rect 22340 24452 22396 24508
rect 22396 24452 22400 24508
rect 22336 24448 22400 24452
rect 22416 24508 22480 24512
rect 22416 24452 22420 24508
rect 22420 24452 22476 24508
rect 22476 24452 22480 24508
rect 22416 24448 22480 24452
rect 22496 24508 22560 24512
rect 22496 24452 22500 24508
rect 22500 24452 22556 24508
rect 22556 24452 22560 24508
rect 22496 24448 22560 24452
rect 28176 24508 28240 24512
rect 28176 24452 28180 24508
rect 28180 24452 28236 24508
rect 28236 24452 28240 24508
rect 28176 24448 28240 24452
rect 28256 24508 28320 24512
rect 28256 24452 28260 24508
rect 28260 24452 28316 24508
rect 28316 24452 28320 24508
rect 28256 24448 28320 24452
rect 28336 24508 28400 24512
rect 28336 24452 28340 24508
rect 28340 24452 28396 24508
rect 28396 24452 28400 24508
rect 28336 24448 28400 24452
rect 28416 24508 28480 24512
rect 28416 24452 28420 24508
rect 28420 24452 28476 24508
rect 28476 24452 28480 24508
rect 28416 24448 28480 24452
rect 28496 24508 28560 24512
rect 28496 24452 28500 24508
rect 28500 24452 28556 24508
rect 28556 24452 28560 24508
rect 28496 24448 28560 24452
rect 4916 23964 4980 23968
rect 4916 23908 4920 23964
rect 4920 23908 4976 23964
rect 4976 23908 4980 23964
rect 4916 23904 4980 23908
rect 4996 23964 5060 23968
rect 4996 23908 5000 23964
rect 5000 23908 5056 23964
rect 5056 23908 5060 23964
rect 4996 23904 5060 23908
rect 5076 23964 5140 23968
rect 5076 23908 5080 23964
rect 5080 23908 5136 23964
rect 5136 23908 5140 23964
rect 5076 23904 5140 23908
rect 5156 23964 5220 23968
rect 5156 23908 5160 23964
rect 5160 23908 5216 23964
rect 5216 23908 5220 23964
rect 5156 23904 5220 23908
rect 5236 23964 5300 23968
rect 5236 23908 5240 23964
rect 5240 23908 5296 23964
rect 5296 23908 5300 23964
rect 5236 23904 5300 23908
rect 10916 23964 10980 23968
rect 10916 23908 10920 23964
rect 10920 23908 10976 23964
rect 10976 23908 10980 23964
rect 10916 23904 10980 23908
rect 10996 23964 11060 23968
rect 10996 23908 11000 23964
rect 11000 23908 11056 23964
rect 11056 23908 11060 23964
rect 10996 23904 11060 23908
rect 11076 23964 11140 23968
rect 11076 23908 11080 23964
rect 11080 23908 11136 23964
rect 11136 23908 11140 23964
rect 11076 23904 11140 23908
rect 11156 23964 11220 23968
rect 11156 23908 11160 23964
rect 11160 23908 11216 23964
rect 11216 23908 11220 23964
rect 11156 23904 11220 23908
rect 11236 23964 11300 23968
rect 11236 23908 11240 23964
rect 11240 23908 11296 23964
rect 11296 23908 11300 23964
rect 11236 23904 11300 23908
rect 16916 23964 16980 23968
rect 16916 23908 16920 23964
rect 16920 23908 16976 23964
rect 16976 23908 16980 23964
rect 16916 23904 16980 23908
rect 16996 23964 17060 23968
rect 16996 23908 17000 23964
rect 17000 23908 17056 23964
rect 17056 23908 17060 23964
rect 16996 23904 17060 23908
rect 17076 23964 17140 23968
rect 17076 23908 17080 23964
rect 17080 23908 17136 23964
rect 17136 23908 17140 23964
rect 17076 23904 17140 23908
rect 17156 23964 17220 23968
rect 17156 23908 17160 23964
rect 17160 23908 17216 23964
rect 17216 23908 17220 23964
rect 17156 23904 17220 23908
rect 17236 23964 17300 23968
rect 17236 23908 17240 23964
rect 17240 23908 17296 23964
rect 17296 23908 17300 23964
rect 17236 23904 17300 23908
rect 22916 23964 22980 23968
rect 22916 23908 22920 23964
rect 22920 23908 22976 23964
rect 22976 23908 22980 23964
rect 22916 23904 22980 23908
rect 22996 23964 23060 23968
rect 22996 23908 23000 23964
rect 23000 23908 23056 23964
rect 23056 23908 23060 23964
rect 22996 23904 23060 23908
rect 23076 23964 23140 23968
rect 23076 23908 23080 23964
rect 23080 23908 23136 23964
rect 23136 23908 23140 23964
rect 23076 23904 23140 23908
rect 23156 23964 23220 23968
rect 23156 23908 23160 23964
rect 23160 23908 23216 23964
rect 23216 23908 23220 23964
rect 23156 23904 23220 23908
rect 23236 23964 23300 23968
rect 23236 23908 23240 23964
rect 23240 23908 23296 23964
rect 23296 23908 23300 23964
rect 23236 23904 23300 23908
rect 28916 23964 28980 23968
rect 28916 23908 28920 23964
rect 28920 23908 28976 23964
rect 28976 23908 28980 23964
rect 28916 23904 28980 23908
rect 28996 23964 29060 23968
rect 28996 23908 29000 23964
rect 29000 23908 29056 23964
rect 29056 23908 29060 23964
rect 28996 23904 29060 23908
rect 29076 23964 29140 23968
rect 29076 23908 29080 23964
rect 29080 23908 29136 23964
rect 29136 23908 29140 23964
rect 29076 23904 29140 23908
rect 29156 23964 29220 23968
rect 29156 23908 29160 23964
rect 29160 23908 29216 23964
rect 29216 23908 29220 23964
rect 29156 23904 29220 23908
rect 29236 23964 29300 23968
rect 29236 23908 29240 23964
rect 29240 23908 29296 23964
rect 29296 23908 29300 23964
rect 29236 23904 29300 23908
rect 14228 23428 14292 23492
rect 4176 23420 4240 23424
rect 4176 23364 4180 23420
rect 4180 23364 4236 23420
rect 4236 23364 4240 23420
rect 4176 23360 4240 23364
rect 4256 23420 4320 23424
rect 4256 23364 4260 23420
rect 4260 23364 4316 23420
rect 4316 23364 4320 23420
rect 4256 23360 4320 23364
rect 4336 23420 4400 23424
rect 4336 23364 4340 23420
rect 4340 23364 4396 23420
rect 4396 23364 4400 23420
rect 4336 23360 4400 23364
rect 4416 23420 4480 23424
rect 4416 23364 4420 23420
rect 4420 23364 4476 23420
rect 4476 23364 4480 23420
rect 4416 23360 4480 23364
rect 4496 23420 4560 23424
rect 4496 23364 4500 23420
rect 4500 23364 4556 23420
rect 4556 23364 4560 23420
rect 4496 23360 4560 23364
rect 10176 23420 10240 23424
rect 10176 23364 10180 23420
rect 10180 23364 10236 23420
rect 10236 23364 10240 23420
rect 10176 23360 10240 23364
rect 10256 23420 10320 23424
rect 10256 23364 10260 23420
rect 10260 23364 10316 23420
rect 10316 23364 10320 23420
rect 10256 23360 10320 23364
rect 10336 23420 10400 23424
rect 10336 23364 10340 23420
rect 10340 23364 10396 23420
rect 10396 23364 10400 23420
rect 10336 23360 10400 23364
rect 10416 23420 10480 23424
rect 10416 23364 10420 23420
rect 10420 23364 10476 23420
rect 10476 23364 10480 23420
rect 10416 23360 10480 23364
rect 10496 23420 10560 23424
rect 10496 23364 10500 23420
rect 10500 23364 10556 23420
rect 10556 23364 10560 23420
rect 10496 23360 10560 23364
rect 16176 23420 16240 23424
rect 16176 23364 16180 23420
rect 16180 23364 16236 23420
rect 16236 23364 16240 23420
rect 16176 23360 16240 23364
rect 16256 23420 16320 23424
rect 16256 23364 16260 23420
rect 16260 23364 16316 23420
rect 16316 23364 16320 23420
rect 16256 23360 16320 23364
rect 16336 23420 16400 23424
rect 16336 23364 16340 23420
rect 16340 23364 16396 23420
rect 16396 23364 16400 23420
rect 16336 23360 16400 23364
rect 16416 23420 16480 23424
rect 16416 23364 16420 23420
rect 16420 23364 16476 23420
rect 16476 23364 16480 23420
rect 16416 23360 16480 23364
rect 16496 23420 16560 23424
rect 16496 23364 16500 23420
rect 16500 23364 16556 23420
rect 16556 23364 16560 23420
rect 16496 23360 16560 23364
rect 22176 23420 22240 23424
rect 22176 23364 22180 23420
rect 22180 23364 22236 23420
rect 22236 23364 22240 23420
rect 22176 23360 22240 23364
rect 22256 23420 22320 23424
rect 22256 23364 22260 23420
rect 22260 23364 22316 23420
rect 22316 23364 22320 23420
rect 22256 23360 22320 23364
rect 22336 23420 22400 23424
rect 22336 23364 22340 23420
rect 22340 23364 22396 23420
rect 22396 23364 22400 23420
rect 22336 23360 22400 23364
rect 22416 23420 22480 23424
rect 22416 23364 22420 23420
rect 22420 23364 22476 23420
rect 22476 23364 22480 23420
rect 22416 23360 22480 23364
rect 22496 23420 22560 23424
rect 22496 23364 22500 23420
rect 22500 23364 22556 23420
rect 22556 23364 22560 23420
rect 22496 23360 22560 23364
rect 28176 23420 28240 23424
rect 28176 23364 28180 23420
rect 28180 23364 28236 23420
rect 28236 23364 28240 23420
rect 28176 23360 28240 23364
rect 28256 23420 28320 23424
rect 28256 23364 28260 23420
rect 28260 23364 28316 23420
rect 28316 23364 28320 23420
rect 28256 23360 28320 23364
rect 28336 23420 28400 23424
rect 28336 23364 28340 23420
rect 28340 23364 28396 23420
rect 28396 23364 28400 23420
rect 28336 23360 28400 23364
rect 28416 23420 28480 23424
rect 28416 23364 28420 23420
rect 28420 23364 28476 23420
rect 28476 23364 28480 23420
rect 28416 23360 28480 23364
rect 28496 23420 28560 23424
rect 28496 23364 28500 23420
rect 28500 23364 28556 23420
rect 28556 23364 28560 23420
rect 28496 23360 28560 23364
rect 4916 22876 4980 22880
rect 4916 22820 4920 22876
rect 4920 22820 4976 22876
rect 4976 22820 4980 22876
rect 4916 22816 4980 22820
rect 4996 22876 5060 22880
rect 4996 22820 5000 22876
rect 5000 22820 5056 22876
rect 5056 22820 5060 22876
rect 4996 22816 5060 22820
rect 5076 22876 5140 22880
rect 5076 22820 5080 22876
rect 5080 22820 5136 22876
rect 5136 22820 5140 22876
rect 5076 22816 5140 22820
rect 5156 22876 5220 22880
rect 5156 22820 5160 22876
rect 5160 22820 5216 22876
rect 5216 22820 5220 22876
rect 5156 22816 5220 22820
rect 5236 22876 5300 22880
rect 5236 22820 5240 22876
rect 5240 22820 5296 22876
rect 5296 22820 5300 22876
rect 5236 22816 5300 22820
rect 10916 22876 10980 22880
rect 10916 22820 10920 22876
rect 10920 22820 10976 22876
rect 10976 22820 10980 22876
rect 10916 22816 10980 22820
rect 10996 22876 11060 22880
rect 10996 22820 11000 22876
rect 11000 22820 11056 22876
rect 11056 22820 11060 22876
rect 10996 22816 11060 22820
rect 11076 22876 11140 22880
rect 11076 22820 11080 22876
rect 11080 22820 11136 22876
rect 11136 22820 11140 22876
rect 11076 22816 11140 22820
rect 11156 22876 11220 22880
rect 11156 22820 11160 22876
rect 11160 22820 11216 22876
rect 11216 22820 11220 22876
rect 11156 22816 11220 22820
rect 11236 22876 11300 22880
rect 11236 22820 11240 22876
rect 11240 22820 11296 22876
rect 11296 22820 11300 22876
rect 11236 22816 11300 22820
rect 16916 22876 16980 22880
rect 16916 22820 16920 22876
rect 16920 22820 16976 22876
rect 16976 22820 16980 22876
rect 16916 22816 16980 22820
rect 16996 22876 17060 22880
rect 16996 22820 17000 22876
rect 17000 22820 17056 22876
rect 17056 22820 17060 22876
rect 16996 22816 17060 22820
rect 17076 22876 17140 22880
rect 17076 22820 17080 22876
rect 17080 22820 17136 22876
rect 17136 22820 17140 22876
rect 17076 22816 17140 22820
rect 17156 22876 17220 22880
rect 17156 22820 17160 22876
rect 17160 22820 17216 22876
rect 17216 22820 17220 22876
rect 17156 22816 17220 22820
rect 17236 22876 17300 22880
rect 17236 22820 17240 22876
rect 17240 22820 17296 22876
rect 17296 22820 17300 22876
rect 17236 22816 17300 22820
rect 22916 22876 22980 22880
rect 22916 22820 22920 22876
rect 22920 22820 22976 22876
rect 22976 22820 22980 22876
rect 22916 22816 22980 22820
rect 22996 22876 23060 22880
rect 22996 22820 23000 22876
rect 23000 22820 23056 22876
rect 23056 22820 23060 22876
rect 22996 22816 23060 22820
rect 23076 22876 23140 22880
rect 23076 22820 23080 22876
rect 23080 22820 23136 22876
rect 23136 22820 23140 22876
rect 23076 22816 23140 22820
rect 23156 22876 23220 22880
rect 23156 22820 23160 22876
rect 23160 22820 23216 22876
rect 23216 22820 23220 22876
rect 23156 22816 23220 22820
rect 23236 22876 23300 22880
rect 23236 22820 23240 22876
rect 23240 22820 23296 22876
rect 23296 22820 23300 22876
rect 23236 22816 23300 22820
rect 28916 22876 28980 22880
rect 28916 22820 28920 22876
rect 28920 22820 28976 22876
rect 28976 22820 28980 22876
rect 28916 22816 28980 22820
rect 28996 22876 29060 22880
rect 28996 22820 29000 22876
rect 29000 22820 29056 22876
rect 29056 22820 29060 22876
rect 28996 22816 29060 22820
rect 29076 22876 29140 22880
rect 29076 22820 29080 22876
rect 29080 22820 29136 22876
rect 29136 22820 29140 22876
rect 29076 22816 29140 22820
rect 29156 22876 29220 22880
rect 29156 22820 29160 22876
rect 29160 22820 29216 22876
rect 29216 22820 29220 22876
rect 29156 22816 29220 22820
rect 29236 22876 29300 22880
rect 29236 22820 29240 22876
rect 29240 22820 29296 22876
rect 29296 22820 29300 22876
rect 29236 22816 29300 22820
rect 4176 22332 4240 22336
rect 4176 22276 4180 22332
rect 4180 22276 4236 22332
rect 4236 22276 4240 22332
rect 4176 22272 4240 22276
rect 4256 22332 4320 22336
rect 4256 22276 4260 22332
rect 4260 22276 4316 22332
rect 4316 22276 4320 22332
rect 4256 22272 4320 22276
rect 4336 22332 4400 22336
rect 4336 22276 4340 22332
rect 4340 22276 4396 22332
rect 4396 22276 4400 22332
rect 4336 22272 4400 22276
rect 4416 22332 4480 22336
rect 4416 22276 4420 22332
rect 4420 22276 4476 22332
rect 4476 22276 4480 22332
rect 4416 22272 4480 22276
rect 4496 22332 4560 22336
rect 4496 22276 4500 22332
rect 4500 22276 4556 22332
rect 4556 22276 4560 22332
rect 4496 22272 4560 22276
rect 10176 22332 10240 22336
rect 10176 22276 10180 22332
rect 10180 22276 10236 22332
rect 10236 22276 10240 22332
rect 10176 22272 10240 22276
rect 10256 22332 10320 22336
rect 10256 22276 10260 22332
rect 10260 22276 10316 22332
rect 10316 22276 10320 22332
rect 10256 22272 10320 22276
rect 10336 22332 10400 22336
rect 10336 22276 10340 22332
rect 10340 22276 10396 22332
rect 10396 22276 10400 22332
rect 10336 22272 10400 22276
rect 10416 22332 10480 22336
rect 10416 22276 10420 22332
rect 10420 22276 10476 22332
rect 10476 22276 10480 22332
rect 10416 22272 10480 22276
rect 10496 22332 10560 22336
rect 10496 22276 10500 22332
rect 10500 22276 10556 22332
rect 10556 22276 10560 22332
rect 10496 22272 10560 22276
rect 16176 22332 16240 22336
rect 16176 22276 16180 22332
rect 16180 22276 16236 22332
rect 16236 22276 16240 22332
rect 16176 22272 16240 22276
rect 16256 22332 16320 22336
rect 16256 22276 16260 22332
rect 16260 22276 16316 22332
rect 16316 22276 16320 22332
rect 16256 22272 16320 22276
rect 16336 22332 16400 22336
rect 16336 22276 16340 22332
rect 16340 22276 16396 22332
rect 16396 22276 16400 22332
rect 16336 22272 16400 22276
rect 16416 22332 16480 22336
rect 16416 22276 16420 22332
rect 16420 22276 16476 22332
rect 16476 22276 16480 22332
rect 16416 22272 16480 22276
rect 16496 22332 16560 22336
rect 16496 22276 16500 22332
rect 16500 22276 16556 22332
rect 16556 22276 16560 22332
rect 16496 22272 16560 22276
rect 22176 22332 22240 22336
rect 22176 22276 22180 22332
rect 22180 22276 22236 22332
rect 22236 22276 22240 22332
rect 22176 22272 22240 22276
rect 22256 22332 22320 22336
rect 22256 22276 22260 22332
rect 22260 22276 22316 22332
rect 22316 22276 22320 22332
rect 22256 22272 22320 22276
rect 22336 22332 22400 22336
rect 22336 22276 22340 22332
rect 22340 22276 22396 22332
rect 22396 22276 22400 22332
rect 22336 22272 22400 22276
rect 22416 22332 22480 22336
rect 22416 22276 22420 22332
rect 22420 22276 22476 22332
rect 22476 22276 22480 22332
rect 22416 22272 22480 22276
rect 22496 22332 22560 22336
rect 22496 22276 22500 22332
rect 22500 22276 22556 22332
rect 22556 22276 22560 22332
rect 22496 22272 22560 22276
rect 28176 22332 28240 22336
rect 28176 22276 28180 22332
rect 28180 22276 28236 22332
rect 28236 22276 28240 22332
rect 28176 22272 28240 22276
rect 28256 22332 28320 22336
rect 28256 22276 28260 22332
rect 28260 22276 28316 22332
rect 28316 22276 28320 22332
rect 28256 22272 28320 22276
rect 28336 22332 28400 22336
rect 28336 22276 28340 22332
rect 28340 22276 28396 22332
rect 28396 22276 28400 22332
rect 28336 22272 28400 22276
rect 28416 22332 28480 22336
rect 28416 22276 28420 22332
rect 28420 22276 28476 22332
rect 28476 22276 28480 22332
rect 28416 22272 28480 22276
rect 28496 22332 28560 22336
rect 28496 22276 28500 22332
rect 28500 22276 28556 22332
rect 28556 22276 28560 22332
rect 28496 22272 28560 22276
rect 4916 21788 4980 21792
rect 4916 21732 4920 21788
rect 4920 21732 4976 21788
rect 4976 21732 4980 21788
rect 4916 21728 4980 21732
rect 4996 21788 5060 21792
rect 4996 21732 5000 21788
rect 5000 21732 5056 21788
rect 5056 21732 5060 21788
rect 4996 21728 5060 21732
rect 5076 21788 5140 21792
rect 5076 21732 5080 21788
rect 5080 21732 5136 21788
rect 5136 21732 5140 21788
rect 5076 21728 5140 21732
rect 5156 21788 5220 21792
rect 5156 21732 5160 21788
rect 5160 21732 5216 21788
rect 5216 21732 5220 21788
rect 5156 21728 5220 21732
rect 5236 21788 5300 21792
rect 5236 21732 5240 21788
rect 5240 21732 5296 21788
rect 5296 21732 5300 21788
rect 5236 21728 5300 21732
rect 10916 21788 10980 21792
rect 10916 21732 10920 21788
rect 10920 21732 10976 21788
rect 10976 21732 10980 21788
rect 10916 21728 10980 21732
rect 10996 21788 11060 21792
rect 10996 21732 11000 21788
rect 11000 21732 11056 21788
rect 11056 21732 11060 21788
rect 10996 21728 11060 21732
rect 11076 21788 11140 21792
rect 11076 21732 11080 21788
rect 11080 21732 11136 21788
rect 11136 21732 11140 21788
rect 11076 21728 11140 21732
rect 11156 21788 11220 21792
rect 11156 21732 11160 21788
rect 11160 21732 11216 21788
rect 11216 21732 11220 21788
rect 11156 21728 11220 21732
rect 11236 21788 11300 21792
rect 11236 21732 11240 21788
rect 11240 21732 11296 21788
rect 11296 21732 11300 21788
rect 11236 21728 11300 21732
rect 16916 21788 16980 21792
rect 16916 21732 16920 21788
rect 16920 21732 16976 21788
rect 16976 21732 16980 21788
rect 16916 21728 16980 21732
rect 16996 21788 17060 21792
rect 16996 21732 17000 21788
rect 17000 21732 17056 21788
rect 17056 21732 17060 21788
rect 16996 21728 17060 21732
rect 17076 21788 17140 21792
rect 17076 21732 17080 21788
rect 17080 21732 17136 21788
rect 17136 21732 17140 21788
rect 17076 21728 17140 21732
rect 17156 21788 17220 21792
rect 17156 21732 17160 21788
rect 17160 21732 17216 21788
rect 17216 21732 17220 21788
rect 17156 21728 17220 21732
rect 17236 21788 17300 21792
rect 17236 21732 17240 21788
rect 17240 21732 17296 21788
rect 17296 21732 17300 21788
rect 17236 21728 17300 21732
rect 22916 21788 22980 21792
rect 22916 21732 22920 21788
rect 22920 21732 22976 21788
rect 22976 21732 22980 21788
rect 22916 21728 22980 21732
rect 22996 21788 23060 21792
rect 22996 21732 23000 21788
rect 23000 21732 23056 21788
rect 23056 21732 23060 21788
rect 22996 21728 23060 21732
rect 23076 21788 23140 21792
rect 23076 21732 23080 21788
rect 23080 21732 23136 21788
rect 23136 21732 23140 21788
rect 23076 21728 23140 21732
rect 23156 21788 23220 21792
rect 23156 21732 23160 21788
rect 23160 21732 23216 21788
rect 23216 21732 23220 21788
rect 23156 21728 23220 21732
rect 23236 21788 23300 21792
rect 23236 21732 23240 21788
rect 23240 21732 23296 21788
rect 23296 21732 23300 21788
rect 23236 21728 23300 21732
rect 28916 21788 28980 21792
rect 28916 21732 28920 21788
rect 28920 21732 28976 21788
rect 28976 21732 28980 21788
rect 28916 21728 28980 21732
rect 28996 21788 29060 21792
rect 28996 21732 29000 21788
rect 29000 21732 29056 21788
rect 29056 21732 29060 21788
rect 28996 21728 29060 21732
rect 29076 21788 29140 21792
rect 29076 21732 29080 21788
rect 29080 21732 29136 21788
rect 29136 21732 29140 21788
rect 29076 21728 29140 21732
rect 29156 21788 29220 21792
rect 29156 21732 29160 21788
rect 29160 21732 29216 21788
rect 29216 21732 29220 21788
rect 29156 21728 29220 21732
rect 29236 21788 29300 21792
rect 29236 21732 29240 21788
rect 29240 21732 29296 21788
rect 29296 21732 29300 21788
rect 29236 21728 29300 21732
rect 4176 21244 4240 21248
rect 4176 21188 4180 21244
rect 4180 21188 4236 21244
rect 4236 21188 4240 21244
rect 4176 21184 4240 21188
rect 4256 21244 4320 21248
rect 4256 21188 4260 21244
rect 4260 21188 4316 21244
rect 4316 21188 4320 21244
rect 4256 21184 4320 21188
rect 4336 21244 4400 21248
rect 4336 21188 4340 21244
rect 4340 21188 4396 21244
rect 4396 21188 4400 21244
rect 4336 21184 4400 21188
rect 4416 21244 4480 21248
rect 4416 21188 4420 21244
rect 4420 21188 4476 21244
rect 4476 21188 4480 21244
rect 4416 21184 4480 21188
rect 4496 21244 4560 21248
rect 4496 21188 4500 21244
rect 4500 21188 4556 21244
rect 4556 21188 4560 21244
rect 4496 21184 4560 21188
rect 10176 21244 10240 21248
rect 10176 21188 10180 21244
rect 10180 21188 10236 21244
rect 10236 21188 10240 21244
rect 10176 21184 10240 21188
rect 10256 21244 10320 21248
rect 10256 21188 10260 21244
rect 10260 21188 10316 21244
rect 10316 21188 10320 21244
rect 10256 21184 10320 21188
rect 10336 21244 10400 21248
rect 10336 21188 10340 21244
rect 10340 21188 10396 21244
rect 10396 21188 10400 21244
rect 10336 21184 10400 21188
rect 10416 21244 10480 21248
rect 10416 21188 10420 21244
rect 10420 21188 10476 21244
rect 10476 21188 10480 21244
rect 10416 21184 10480 21188
rect 10496 21244 10560 21248
rect 10496 21188 10500 21244
rect 10500 21188 10556 21244
rect 10556 21188 10560 21244
rect 10496 21184 10560 21188
rect 16176 21244 16240 21248
rect 16176 21188 16180 21244
rect 16180 21188 16236 21244
rect 16236 21188 16240 21244
rect 16176 21184 16240 21188
rect 16256 21244 16320 21248
rect 16256 21188 16260 21244
rect 16260 21188 16316 21244
rect 16316 21188 16320 21244
rect 16256 21184 16320 21188
rect 16336 21244 16400 21248
rect 16336 21188 16340 21244
rect 16340 21188 16396 21244
rect 16396 21188 16400 21244
rect 16336 21184 16400 21188
rect 16416 21244 16480 21248
rect 16416 21188 16420 21244
rect 16420 21188 16476 21244
rect 16476 21188 16480 21244
rect 16416 21184 16480 21188
rect 16496 21244 16560 21248
rect 16496 21188 16500 21244
rect 16500 21188 16556 21244
rect 16556 21188 16560 21244
rect 16496 21184 16560 21188
rect 22176 21244 22240 21248
rect 22176 21188 22180 21244
rect 22180 21188 22236 21244
rect 22236 21188 22240 21244
rect 22176 21184 22240 21188
rect 22256 21244 22320 21248
rect 22256 21188 22260 21244
rect 22260 21188 22316 21244
rect 22316 21188 22320 21244
rect 22256 21184 22320 21188
rect 22336 21244 22400 21248
rect 22336 21188 22340 21244
rect 22340 21188 22396 21244
rect 22396 21188 22400 21244
rect 22336 21184 22400 21188
rect 22416 21244 22480 21248
rect 22416 21188 22420 21244
rect 22420 21188 22476 21244
rect 22476 21188 22480 21244
rect 22416 21184 22480 21188
rect 22496 21244 22560 21248
rect 22496 21188 22500 21244
rect 22500 21188 22556 21244
rect 22556 21188 22560 21244
rect 22496 21184 22560 21188
rect 28176 21244 28240 21248
rect 28176 21188 28180 21244
rect 28180 21188 28236 21244
rect 28236 21188 28240 21244
rect 28176 21184 28240 21188
rect 28256 21244 28320 21248
rect 28256 21188 28260 21244
rect 28260 21188 28316 21244
rect 28316 21188 28320 21244
rect 28256 21184 28320 21188
rect 28336 21244 28400 21248
rect 28336 21188 28340 21244
rect 28340 21188 28396 21244
rect 28396 21188 28400 21244
rect 28336 21184 28400 21188
rect 28416 21244 28480 21248
rect 28416 21188 28420 21244
rect 28420 21188 28476 21244
rect 28476 21188 28480 21244
rect 28416 21184 28480 21188
rect 28496 21244 28560 21248
rect 28496 21188 28500 21244
rect 28500 21188 28556 21244
rect 28556 21188 28560 21244
rect 28496 21184 28560 21188
rect 12940 20708 13004 20772
rect 20668 20768 20732 20772
rect 20668 20712 20718 20768
rect 20718 20712 20732 20768
rect 20668 20708 20732 20712
rect 4916 20700 4980 20704
rect 4916 20644 4920 20700
rect 4920 20644 4976 20700
rect 4976 20644 4980 20700
rect 4916 20640 4980 20644
rect 4996 20700 5060 20704
rect 4996 20644 5000 20700
rect 5000 20644 5056 20700
rect 5056 20644 5060 20700
rect 4996 20640 5060 20644
rect 5076 20700 5140 20704
rect 5076 20644 5080 20700
rect 5080 20644 5136 20700
rect 5136 20644 5140 20700
rect 5076 20640 5140 20644
rect 5156 20700 5220 20704
rect 5156 20644 5160 20700
rect 5160 20644 5216 20700
rect 5216 20644 5220 20700
rect 5156 20640 5220 20644
rect 5236 20700 5300 20704
rect 5236 20644 5240 20700
rect 5240 20644 5296 20700
rect 5296 20644 5300 20700
rect 5236 20640 5300 20644
rect 10916 20700 10980 20704
rect 10916 20644 10920 20700
rect 10920 20644 10976 20700
rect 10976 20644 10980 20700
rect 10916 20640 10980 20644
rect 10996 20700 11060 20704
rect 10996 20644 11000 20700
rect 11000 20644 11056 20700
rect 11056 20644 11060 20700
rect 10996 20640 11060 20644
rect 11076 20700 11140 20704
rect 11076 20644 11080 20700
rect 11080 20644 11136 20700
rect 11136 20644 11140 20700
rect 11076 20640 11140 20644
rect 11156 20700 11220 20704
rect 11156 20644 11160 20700
rect 11160 20644 11216 20700
rect 11216 20644 11220 20700
rect 11156 20640 11220 20644
rect 11236 20700 11300 20704
rect 11236 20644 11240 20700
rect 11240 20644 11296 20700
rect 11296 20644 11300 20700
rect 11236 20640 11300 20644
rect 16916 20700 16980 20704
rect 16916 20644 16920 20700
rect 16920 20644 16976 20700
rect 16976 20644 16980 20700
rect 16916 20640 16980 20644
rect 16996 20700 17060 20704
rect 16996 20644 17000 20700
rect 17000 20644 17056 20700
rect 17056 20644 17060 20700
rect 16996 20640 17060 20644
rect 17076 20700 17140 20704
rect 17076 20644 17080 20700
rect 17080 20644 17136 20700
rect 17136 20644 17140 20700
rect 17076 20640 17140 20644
rect 17156 20700 17220 20704
rect 17156 20644 17160 20700
rect 17160 20644 17216 20700
rect 17216 20644 17220 20700
rect 17156 20640 17220 20644
rect 17236 20700 17300 20704
rect 17236 20644 17240 20700
rect 17240 20644 17296 20700
rect 17296 20644 17300 20700
rect 17236 20640 17300 20644
rect 22916 20700 22980 20704
rect 22916 20644 22920 20700
rect 22920 20644 22976 20700
rect 22976 20644 22980 20700
rect 22916 20640 22980 20644
rect 22996 20700 23060 20704
rect 22996 20644 23000 20700
rect 23000 20644 23056 20700
rect 23056 20644 23060 20700
rect 22996 20640 23060 20644
rect 23076 20700 23140 20704
rect 23076 20644 23080 20700
rect 23080 20644 23136 20700
rect 23136 20644 23140 20700
rect 23076 20640 23140 20644
rect 23156 20700 23220 20704
rect 23156 20644 23160 20700
rect 23160 20644 23216 20700
rect 23216 20644 23220 20700
rect 23156 20640 23220 20644
rect 23236 20700 23300 20704
rect 23236 20644 23240 20700
rect 23240 20644 23296 20700
rect 23296 20644 23300 20700
rect 23236 20640 23300 20644
rect 28916 20700 28980 20704
rect 28916 20644 28920 20700
rect 28920 20644 28976 20700
rect 28976 20644 28980 20700
rect 28916 20640 28980 20644
rect 28996 20700 29060 20704
rect 28996 20644 29000 20700
rect 29000 20644 29056 20700
rect 29056 20644 29060 20700
rect 28996 20640 29060 20644
rect 29076 20700 29140 20704
rect 29076 20644 29080 20700
rect 29080 20644 29136 20700
rect 29136 20644 29140 20700
rect 29076 20640 29140 20644
rect 29156 20700 29220 20704
rect 29156 20644 29160 20700
rect 29160 20644 29216 20700
rect 29216 20644 29220 20700
rect 29156 20640 29220 20644
rect 29236 20700 29300 20704
rect 29236 20644 29240 20700
rect 29240 20644 29296 20700
rect 29296 20644 29300 20700
rect 29236 20640 29300 20644
rect 4176 20156 4240 20160
rect 4176 20100 4180 20156
rect 4180 20100 4236 20156
rect 4236 20100 4240 20156
rect 4176 20096 4240 20100
rect 4256 20156 4320 20160
rect 4256 20100 4260 20156
rect 4260 20100 4316 20156
rect 4316 20100 4320 20156
rect 4256 20096 4320 20100
rect 4336 20156 4400 20160
rect 4336 20100 4340 20156
rect 4340 20100 4396 20156
rect 4396 20100 4400 20156
rect 4336 20096 4400 20100
rect 4416 20156 4480 20160
rect 4416 20100 4420 20156
rect 4420 20100 4476 20156
rect 4476 20100 4480 20156
rect 4416 20096 4480 20100
rect 4496 20156 4560 20160
rect 4496 20100 4500 20156
rect 4500 20100 4556 20156
rect 4556 20100 4560 20156
rect 4496 20096 4560 20100
rect 10176 20156 10240 20160
rect 10176 20100 10180 20156
rect 10180 20100 10236 20156
rect 10236 20100 10240 20156
rect 10176 20096 10240 20100
rect 10256 20156 10320 20160
rect 10256 20100 10260 20156
rect 10260 20100 10316 20156
rect 10316 20100 10320 20156
rect 10256 20096 10320 20100
rect 10336 20156 10400 20160
rect 10336 20100 10340 20156
rect 10340 20100 10396 20156
rect 10396 20100 10400 20156
rect 10336 20096 10400 20100
rect 10416 20156 10480 20160
rect 10416 20100 10420 20156
rect 10420 20100 10476 20156
rect 10476 20100 10480 20156
rect 10416 20096 10480 20100
rect 10496 20156 10560 20160
rect 10496 20100 10500 20156
rect 10500 20100 10556 20156
rect 10556 20100 10560 20156
rect 10496 20096 10560 20100
rect 16176 20156 16240 20160
rect 16176 20100 16180 20156
rect 16180 20100 16236 20156
rect 16236 20100 16240 20156
rect 16176 20096 16240 20100
rect 16256 20156 16320 20160
rect 16256 20100 16260 20156
rect 16260 20100 16316 20156
rect 16316 20100 16320 20156
rect 16256 20096 16320 20100
rect 16336 20156 16400 20160
rect 16336 20100 16340 20156
rect 16340 20100 16396 20156
rect 16396 20100 16400 20156
rect 16336 20096 16400 20100
rect 16416 20156 16480 20160
rect 16416 20100 16420 20156
rect 16420 20100 16476 20156
rect 16476 20100 16480 20156
rect 16416 20096 16480 20100
rect 16496 20156 16560 20160
rect 16496 20100 16500 20156
rect 16500 20100 16556 20156
rect 16556 20100 16560 20156
rect 16496 20096 16560 20100
rect 22176 20156 22240 20160
rect 22176 20100 22180 20156
rect 22180 20100 22236 20156
rect 22236 20100 22240 20156
rect 22176 20096 22240 20100
rect 22256 20156 22320 20160
rect 22256 20100 22260 20156
rect 22260 20100 22316 20156
rect 22316 20100 22320 20156
rect 22256 20096 22320 20100
rect 22336 20156 22400 20160
rect 22336 20100 22340 20156
rect 22340 20100 22396 20156
rect 22396 20100 22400 20156
rect 22336 20096 22400 20100
rect 22416 20156 22480 20160
rect 22416 20100 22420 20156
rect 22420 20100 22476 20156
rect 22476 20100 22480 20156
rect 22416 20096 22480 20100
rect 22496 20156 22560 20160
rect 22496 20100 22500 20156
rect 22500 20100 22556 20156
rect 22556 20100 22560 20156
rect 22496 20096 22560 20100
rect 28176 20156 28240 20160
rect 28176 20100 28180 20156
rect 28180 20100 28236 20156
rect 28236 20100 28240 20156
rect 28176 20096 28240 20100
rect 28256 20156 28320 20160
rect 28256 20100 28260 20156
rect 28260 20100 28316 20156
rect 28316 20100 28320 20156
rect 28256 20096 28320 20100
rect 28336 20156 28400 20160
rect 28336 20100 28340 20156
rect 28340 20100 28396 20156
rect 28396 20100 28400 20156
rect 28336 20096 28400 20100
rect 28416 20156 28480 20160
rect 28416 20100 28420 20156
rect 28420 20100 28476 20156
rect 28476 20100 28480 20156
rect 28416 20096 28480 20100
rect 28496 20156 28560 20160
rect 28496 20100 28500 20156
rect 28500 20100 28556 20156
rect 28556 20100 28560 20156
rect 28496 20096 28560 20100
rect 4916 19612 4980 19616
rect 4916 19556 4920 19612
rect 4920 19556 4976 19612
rect 4976 19556 4980 19612
rect 4916 19552 4980 19556
rect 4996 19612 5060 19616
rect 4996 19556 5000 19612
rect 5000 19556 5056 19612
rect 5056 19556 5060 19612
rect 4996 19552 5060 19556
rect 5076 19612 5140 19616
rect 5076 19556 5080 19612
rect 5080 19556 5136 19612
rect 5136 19556 5140 19612
rect 5076 19552 5140 19556
rect 5156 19612 5220 19616
rect 5156 19556 5160 19612
rect 5160 19556 5216 19612
rect 5216 19556 5220 19612
rect 5156 19552 5220 19556
rect 5236 19612 5300 19616
rect 5236 19556 5240 19612
rect 5240 19556 5296 19612
rect 5296 19556 5300 19612
rect 5236 19552 5300 19556
rect 10916 19612 10980 19616
rect 10916 19556 10920 19612
rect 10920 19556 10976 19612
rect 10976 19556 10980 19612
rect 10916 19552 10980 19556
rect 10996 19612 11060 19616
rect 10996 19556 11000 19612
rect 11000 19556 11056 19612
rect 11056 19556 11060 19612
rect 10996 19552 11060 19556
rect 11076 19612 11140 19616
rect 11076 19556 11080 19612
rect 11080 19556 11136 19612
rect 11136 19556 11140 19612
rect 11076 19552 11140 19556
rect 11156 19612 11220 19616
rect 11156 19556 11160 19612
rect 11160 19556 11216 19612
rect 11216 19556 11220 19612
rect 11156 19552 11220 19556
rect 11236 19612 11300 19616
rect 11236 19556 11240 19612
rect 11240 19556 11296 19612
rect 11296 19556 11300 19612
rect 11236 19552 11300 19556
rect 16916 19612 16980 19616
rect 16916 19556 16920 19612
rect 16920 19556 16976 19612
rect 16976 19556 16980 19612
rect 16916 19552 16980 19556
rect 16996 19612 17060 19616
rect 16996 19556 17000 19612
rect 17000 19556 17056 19612
rect 17056 19556 17060 19612
rect 16996 19552 17060 19556
rect 17076 19612 17140 19616
rect 17076 19556 17080 19612
rect 17080 19556 17136 19612
rect 17136 19556 17140 19612
rect 17076 19552 17140 19556
rect 17156 19612 17220 19616
rect 17156 19556 17160 19612
rect 17160 19556 17216 19612
rect 17216 19556 17220 19612
rect 17156 19552 17220 19556
rect 17236 19612 17300 19616
rect 17236 19556 17240 19612
rect 17240 19556 17296 19612
rect 17296 19556 17300 19612
rect 17236 19552 17300 19556
rect 22916 19612 22980 19616
rect 22916 19556 22920 19612
rect 22920 19556 22976 19612
rect 22976 19556 22980 19612
rect 22916 19552 22980 19556
rect 22996 19612 23060 19616
rect 22996 19556 23000 19612
rect 23000 19556 23056 19612
rect 23056 19556 23060 19612
rect 22996 19552 23060 19556
rect 23076 19612 23140 19616
rect 23076 19556 23080 19612
rect 23080 19556 23136 19612
rect 23136 19556 23140 19612
rect 23076 19552 23140 19556
rect 23156 19612 23220 19616
rect 23156 19556 23160 19612
rect 23160 19556 23216 19612
rect 23216 19556 23220 19612
rect 23156 19552 23220 19556
rect 23236 19612 23300 19616
rect 23236 19556 23240 19612
rect 23240 19556 23296 19612
rect 23296 19556 23300 19612
rect 23236 19552 23300 19556
rect 28916 19612 28980 19616
rect 28916 19556 28920 19612
rect 28920 19556 28976 19612
rect 28976 19556 28980 19612
rect 28916 19552 28980 19556
rect 28996 19612 29060 19616
rect 28996 19556 29000 19612
rect 29000 19556 29056 19612
rect 29056 19556 29060 19612
rect 28996 19552 29060 19556
rect 29076 19612 29140 19616
rect 29076 19556 29080 19612
rect 29080 19556 29136 19612
rect 29136 19556 29140 19612
rect 29076 19552 29140 19556
rect 29156 19612 29220 19616
rect 29156 19556 29160 19612
rect 29160 19556 29216 19612
rect 29216 19556 29220 19612
rect 29156 19552 29220 19556
rect 29236 19612 29300 19616
rect 29236 19556 29240 19612
rect 29240 19556 29296 19612
rect 29296 19556 29300 19612
rect 29236 19552 29300 19556
rect 14228 19348 14292 19412
rect 4176 19068 4240 19072
rect 4176 19012 4180 19068
rect 4180 19012 4236 19068
rect 4236 19012 4240 19068
rect 4176 19008 4240 19012
rect 4256 19068 4320 19072
rect 4256 19012 4260 19068
rect 4260 19012 4316 19068
rect 4316 19012 4320 19068
rect 4256 19008 4320 19012
rect 4336 19068 4400 19072
rect 4336 19012 4340 19068
rect 4340 19012 4396 19068
rect 4396 19012 4400 19068
rect 4336 19008 4400 19012
rect 4416 19068 4480 19072
rect 4416 19012 4420 19068
rect 4420 19012 4476 19068
rect 4476 19012 4480 19068
rect 4416 19008 4480 19012
rect 4496 19068 4560 19072
rect 4496 19012 4500 19068
rect 4500 19012 4556 19068
rect 4556 19012 4560 19068
rect 4496 19008 4560 19012
rect 10176 19068 10240 19072
rect 10176 19012 10180 19068
rect 10180 19012 10236 19068
rect 10236 19012 10240 19068
rect 10176 19008 10240 19012
rect 10256 19068 10320 19072
rect 10256 19012 10260 19068
rect 10260 19012 10316 19068
rect 10316 19012 10320 19068
rect 10256 19008 10320 19012
rect 10336 19068 10400 19072
rect 10336 19012 10340 19068
rect 10340 19012 10396 19068
rect 10396 19012 10400 19068
rect 10336 19008 10400 19012
rect 10416 19068 10480 19072
rect 10416 19012 10420 19068
rect 10420 19012 10476 19068
rect 10476 19012 10480 19068
rect 10416 19008 10480 19012
rect 10496 19068 10560 19072
rect 10496 19012 10500 19068
rect 10500 19012 10556 19068
rect 10556 19012 10560 19068
rect 10496 19008 10560 19012
rect 16176 19068 16240 19072
rect 16176 19012 16180 19068
rect 16180 19012 16236 19068
rect 16236 19012 16240 19068
rect 16176 19008 16240 19012
rect 16256 19068 16320 19072
rect 16256 19012 16260 19068
rect 16260 19012 16316 19068
rect 16316 19012 16320 19068
rect 16256 19008 16320 19012
rect 16336 19068 16400 19072
rect 16336 19012 16340 19068
rect 16340 19012 16396 19068
rect 16396 19012 16400 19068
rect 16336 19008 16400 19012
rect 16416 19068 16480 19072
rect 16416 19012 16420 19068
rect 16420 19012 16476 19068
rect 16476 19012 16480 19068
rect 16416 19008 16480 19012
rect 16496 19068 16560 19072
rect 16496 19012 16500 19068
rect 16500 19012 16556 19068
rect 16556 19012 16560 19068
rect 16496 19008 16560 19012
rect 22176 19068 22240 19072
rect 22176 19012 22180 19068
rect 22180 19012 22236 19068
rect 22236 19012 22240 19068
rect 22176 19008 22240 19012
rect 22256 19068 22320 19072
rect 22256 19012 22260 19068
rect 22260 19012 22316 19068
rect 22316 19012 22320 19068
rect 22256 19008 22320 19012
rect 22336 19068 22400 19072
rect 22336 19012 22340 19068
rect 22340 19012 22396 19068
rect 22396 19012 22400 19068
rect 22336 19008 22400 19012
rect 22416 19068 22480 19072
rect 22416 19012 22420 19068
rect 22420 19012 22476 19068
rect 22476 19012 22480 19068
rect 22416 19008 22480 19012
rect 22496 19068 22560 19072
rect 22496 19012 22500 19068
rect 22500 19012 22556 19068
rect 22556 19012 22560 19068
rect 22496 19008 22560 19012
rect 28176 19068 28240 19072
rect 28176 19012 28180 19068
rect 28180 19012 28236 19068
rect 28236 19012 28240 19068
rect 28176 19008 28240 19012
rect 28256 19068 28320 19072
rect 28256 19012 28260 19068
rect 28260 19012 28316 19068
rect 28316 19012 28320 19068
rect 28256 19008 28320 19012
rect 28336 19068 28400 19072
rect 28336 19012 28340 19068
rect 28340 19012 28396 19068
rect 28396 19012 28400 19068
rect 28336 19008 28400 19012
rect 28416 19068 28480 19072
rect 28416 19012 28420 19068
rect 28420 19012 28476 19068
rect 28476 19012 28480 19068
rect 28416 19008 28480 19012
rect 28496 19068 28560 19072
rect 28496 19012 28500 19068
rect 28500 19012 28556 19068
rect 28556 19012 28560 19068
rect 28496 19008 28560 19012
rect 4916 18524 4980 18528
rect 4916 18468 4920 18524
rect 4920 18468 4976 18524
rect 4976 18468 4980 18524
rect 4916 18464 4980 18468
rect 4996 18524 5060 18528
rect 4996 18468 5000 18524
rect 5000 18468 5056 18524
rect 5056 18468 5060 18524
rect 4996 18464 5060 18468
rect 5076 18524 5140 18528
rect 5076 18468 5080 18524
rect 5080 18468 5136 18524
rect 5136 18468 5140 18524
rect 5076 18464 5140 18468
rect 5156 18524 5220 18528
rect 5156 18468 5160 18524
rect 5160 18468 5216 18524
rect 5216 18468 5220 18524
rect 5156 18464 5220 18468
rect 5236 18524 5300 18528
rect 5236 18468 5240 18524
rect 5240 18468 5296 18524
rect 5296 18468 5300 18524
rect 5236 18464 5300 18468
rect 10916 18524 10980 18528
rect 10916 18468 10920 18524
rect 10920 18468 10976 18524
rect 10976 18468 10980 18524
rect 10916 18464 10980 18468
rect 10996 18524 11060 18528
rect 10996 18468 11000 18524
rect 11000 18468 11056 18524
rect 11056 18468 11060 18524
rect 10996 18464 11060 18468
rect 11076 18524 11140 18528
rect 11076 18468 11080 18524
rect 11080 18468 11136 18524
rect 11136 18468 11140 18524
rect 11076 18464 11140 18468
rect 11156 18524 11220 18528
rect 11156 18468 11160 18524
rect 11160 18468 11216 18524
rect 11216 18468 11220 18524
rect 11156 18464 11220 18468
rect 11236 18524 11300 18528
rect 11236 18468 11240 18524
rect 11240 18468 11296 18524
rect 11296 18468 11300 18524
rect 11236 18464 11300 18468
rect 16916 18524 16980 18528
rect 16916 18468 16920 18524
rect 16920 18468 16976 18524
rect 16976 18468 16980 18524
rect 16916 18464 16980 18468
rect 16996 18524 17060 18528
rect 16996 18468 17000 18524
rect 17000 18468 17056 18524
rect 17056 18468 17060 18524
rect 16996 18464 17060 18468
rect 17076 18524 17140 18528
rect 17076 18468 17080 18524
rect 17080 18468 17136 18524
rect 17136 18468 17140 18524
rect 17076 18464 17140 18468
rect 17156 18524 17220 18528
rect 17156 18468 17160 18524
rect 17160 18468 17216 18524
rect 17216 18468 17220 18524
rect 17156 18464 17220 18468
rect 17236 18524 17300 18528
rect 17236 18468 17240 18524
rect 17240 18468 17296 18524
rect 17296 18468 17300 18524
rect 17236 18464 17300 18468
rect 22916 18524 22980 18528
rect 22916 18468 22920 18524
rect 22920 18468 22976 18524
rect 22976 18468 22980 18524
rect 22916 18464 22980 18468
rect 22996 18524 23060 18528
rect 22996 18468 23000 18524
rect 23000 18468 23056 18524
rect 23056 18468 23060 18524
rect 22996 18464 23060 18468
rect 23076 18524 23140 18528
rect 23076 18468 23080 18524
rect 23080 18468 23136 18524
rect 23136 18468 23140 18524
rect 23076 18464 23140 18468
rect 23156 18524 23220 18528
rect 23156 18468 23160 18524
rect 23160 18468 23216 18524
rect 23216 18468 23220 18524
rect 23156 18464 23220 18468
rect 23236 18524 23300 18528
rect 23236 18468 23240 18524
rect 23240 18468 23296 18524
rect 23296 18468 23300 18524
rect 23236 18464 23300 18468
rect 28916 18524 28980 18528
rect 28916 18468 28920 18524
rect 28920 18468 28976 18524
rect 28976 18468 28980 18524
rect 28916 18464 28980 18468
rect 28996 18524 29060 18528
rect 28996 18468 29000 18524
rect 29000 18468 29056 18524
rect 29056 18468 29060 18524
rect 28996 18464 29060 18468
rect 29076 18524 29140 18528
rect 29076 18468 29080 18524
rect 29080 18468 29136 18524
rect 29136 18468 29140 18524
rect 29076 18464 29140 18468
rect 29156 18524 29220 18528
rect 29156 18468 29160 18524
rect 29160 18468 29216 18524
rect 29216 18468 29220 18524
rect 29156 18464 29220 18468
rect 29236 18524 29300 18528
rect 29236 18468 29240 18524
rect 29240 18468 29296 18524
rect 29296 18468 29300 18524
rect 29236 18464 29300 18468
rect 4176 17980 4240 17984
rect 4176 17924 4180 17980
rect 4180 17924 4236 17980
rect 4236 17924 4240 17980
rect 4176 17920 4240 17924
rect 4256 17980 4320 17984
rect 4256 17924 4260 17980
rect 4260 17924 4316 17980
rect 4316 17924 4320 17980
rect 4256 17920 4320 17924
rect 4336 17980 4400 17984
rect 4336 17924 4340 17980
rect 4340 17924 4396 17980
rect 4396 17924 4400 17980
rect 4336 17920 4400 17924
rect 4416 17980 4480 17984
rect 4416 17924 4420 17980
rect 4420 17924 4476 17980
rect 4476 17924 4480 17980
rect 4416 17920 4480 17924
rect 4496 17980 4560 17984
rect 4496 17924 4500 17980
rect 4500 17924 4556 17980
rect 4556 17924 4560 17980
rect 4496 17920 4560 17924
rect 10176 17980 10240 17984
rect 10176 17924 10180 17980
rect 10180 17924 10236 17980
rect 10236 17924 10240 17980
rect 10176 17920 10240 17924
rect 10256 17980 10320 17984
rect 10256 17924 10260 17980
rect 10260 17924 10316 17980
rect 10316 17924 10320 17980
rect 10256 17920 10320 17924
rect 10336 17980 10400 17984
rect 10336 17924 10340 17980
rect 10340 17924 10396 17980
rect 10396 17924 10400 17980
rect 10336 17920 10400 17924
rect 10416 17980 10480 17984
rect 10416 17924 10420 17980
rect 10420 17924 10476 17980
rect 10476 17924 10480 17980
rect 10416 17920 10480 17924
rect 10496 17980 10560 17984
rect 10496 17924 10500 17980
rect 10500 17924 10556 17980
rect 10556 17924 10560 17980
rect 10496 17920 10560 17924
rect 16176 17980 16240 17984
rect 16176 17924 16180 17980
rect 16180 17924 16236 17980
rect 16236 17924 16240 17980
rect 16176 17920 16240 17924
rect 16256 17980 16320 17984
rect 16256 17924 16260 17980
rect 16260 17924 16316 17980
rect 16316 17924 16320 17980
rect 16256 17920 16320 17924
rect 16336 17980 16400 17984
rect 16336 17924 16340 17980
rect 16340 17924 16396 17980
rect 16396 17924 16400 17980
rect 16336 17920 16400 17924
rect 16416 17980 16480 17984
rect 16416 17924 16420 17980
rect 16420 17924 16476 17980
rect 16476 17924 16480 17980
rect 16416 17920 16480 17924
rect 16496 17980 16560 17984
rect 16496 17924 16500 17980
rect 16500 17924 16556 17980
rect 16556 17924 16560 17980
rect 16496 17920 16560 17924
rect 22176 17980 22240 17984
rect 22176 17924 22180 17980
rect 22180 17924 22236 17980
rect 22236 17924 22240 17980
rect 22176 17920 22240 17924
rect 22256 17980 22320 17984
rect 22256 17924 22260 17980
rect 22260 17924 22316 17980
rect 22316 17924 22320 17980
rect 22256 17920 22320 17924
rect 22336 17980 22400 17984
rect 22336 17924 22340 17980
rect 22340 17924 22396 17980
rect 22396 17924 22400 17980
rect 22336 17920 22400 17924
rect 22416 17980 22480 17984
rect 22416 17924 22420 17980
rect 22420 17924 22476 17980
rect 22476 17924 22480 17980
rect 22416 17920 22480 17924
rect 22496 17980 22560 17984
rect 22496 17924 22500 17980
rect 22500 17924 22556 17980
rect 22556 17924 22560 17980
rect 22496 17920 22560 17924
rect 28176 17980 28240 17984
rect 28176 17924 28180 17980
rect 28180 17924 28236 17980
rect 28236 17924 28240 17980
rect 28176 17920 28240 17924
rect 28256 17980 28320 17984
rect 28256 17924 28260 17980
rect 28260 17924 28316 17980
rect 28316 17924 28320 17980
rect 28256 17920 28320 17924
rect 28336 17980 28400 17984
rect 28336 17924 28340 17980
rect 28340 17924 28396 17980
rect 28396 17924 28400 17980
rect 28336 17920 28400 17924
rect 28416 17980 28480 17984
rect 28416 17924 28420 17980
rect 28420 17924 28476 17980
rect 28476 17924 28480 17980
rect 28416 17920 28480 17924
rect 28496 17980 28560 17984
rect 28496 17924 28500 17980
rect 28500 17924 28556 17980
rect 28556 17924 28560 17980
rect 28496 17920 28560 17924
rect 27844 17580 27908 17644
rect 19380 17444 19444 17508
rect 20668 17444 20732 17508
rect 4916 17436 4980 17440
rect 4916 17380 4920 17436
rect 4920 17380 4976 17436
rect 4976 17380 4980 17436
rect 4916 17376 4980 17380
rect 4996 17436 5060 17440
rect 4996 17380 5000 17436
rect 5000 17380 5056 17436
rect 5056 17380 5060 17436
rect 4996 17376 5060 17380
rect 5076 17436 5140 17440
rect 5076 17380 5080 17436
rect 5080 17380 5136 17436
rect 5136 17380 5140 17436
rect 5076 17376 5140 17380
rect 5156 17436 5220 17440
rect 5156 17380 5160 17436
rect 5160 17380 5216 17436
rect 5216 17380 5220 17436
rect 5156 17376 5220 17380
rect 5236 17436 5300 17440
rect 5236 17380 5240 17436
rect 5240 17380 5296 17436
rect 5296 17380 5300 17436
rect 5236 17376 5300 17380
rect 10916 17436 10980 17440
rect 10916 17380 10920 17436
rect 10920 17380 10976 17436
rect 10976 17380 10980 17436
rect 10916 17376 10980 17380
rect 10996 17436 11060 17440
rect 10996 17380 11000 17436
rect 11000 17380 11056 17436
rect 11056 17380 11060 17436
rect 10996 17376 11060 17380
rect 11076 17436 11140 17440
rect 11076 17380 11080 17436
rect 11080 17380 11136 17436
rect 11136 17380 11140 17436
rect 11076 17376 11140 17380
rect 11156 17436 11220 17440
rect 11156 17380 11160 17436
rect 11160 17380 11216 17436
rect 11216 17380 11220 17436
rect 11156 17376 11220 17380
rect 11236 17436 11300 17440
rect 11236 17380 11240 17436
rect 11240 17380 11296 17436
rect 11296 17380 11300 17436
rect 11236 17376 11300 17380
rect 16916 17436 16980 17440
rect 16916 17380 16920 17436
rect 16920 17380 16976 17436
rect 16976 17380 16980 17436
rect 16916 17376 16980 17380
rect 16996 17436 17060 17440
rect 16996 17380 17000 17436
rect 17000 17380 17056 17436
rect 17056 17380 17060 17436
rect 16996 17376 17060 17380
rect 17076 17436 17140 17440
rect 17076 17380 17080 17436
rect 17080 17380 17136 17436
rect 17136 17380 17140 17436
rect 17076 17376 17140 17380
rect 17156 17436 17220 17440
rect 17156 17380 17160 17436
rect 17160 17380 17216 17436
rect 17216 17380 17220 17436
rect 17156 17376 17220 17380
rect 17236 17436 17300 17440
rect 17236 17380 17240 17436
rect 17240 17380 17296 17436
rect 17296 17380 17300 17436
rect 17236 17376 17300 17380
rect 22916 17436 22980 17440
rect 22916 17380 22920 17436
rect 22920 17380 22976 17436
rect 22976 17380 22980 17436
rect 22916 17376 22980 17380
rect 22996 17436 23060 17440
rect 22996 17380 23000 17436
rect 23000 17380 23056 17436
rect 23056 17380 23060 17436
rect 22996 17376 23060 17380
rect 23076 17436 23140 17440
rect 23076 17380 23080 17436
rect 23080 17380 23136 17436
rect 23136 17380 23140 17436
rect 23076 17376 23140 17380
rect 23156 17436 23220 17440
rect 23156 17380 23160 17436
rect 23160 17380 23216 17436
rect 23216 17380 23220 17436
rect 23156 17376 23220 17380
rect 23236 17436 23300 17440
rect 23236 17380 23240 17436
rect 23240 17380 23296 17436
rect 23296 17380 23300 17436
rect 23236 17376 23300 17380
rect 28916 17436 28980 17440
rect 28916 17380 28920 17436
rect 28920 17380 28976 17436
rect 28976 17380 28980 17436
rect 28916 17376 28980 17380
rect 28996 17436 29060 17440
rect 28996 17380 29000 17436
rect 29000 17380 29056 17436
rect 29056 17380 29060 17436
rect 28996 17376 29060 17380
rect 29076 17436 29140 17440
rect 29076 17380 29080 17436
rect 29080 17380 29136 17436
rect 29136 17380 29140 17436
rect 29076 17376 29140 17380
rect 29156 17436 29220 17440
rect 29156 17380 29160 17436
rect 29160 17380 29216 17436
rect 29216 17380 29220 17436
rect 29156 17376 29220 17380
rect 29236 17436 29300 17440
rect 29236 17380 29240 17436
rect 29240 17380 29296 17436
rect 29296 17380 29300 17436
rect 29236 17376 29300 17380
rect 4176 16892 4240 16896
rect 4176 16836 4180 16892
rect 4180 16836 4236 16892
rect 4236 16836 4240 16892
rect 4176 16832 4240 16836
rect 4256 16892 4320 16896
rect 4256 16836 4260 16892
rect 4260 16836 4316 16892
rect 4316 16836 4320 16892
rect 4256 16832 4320 16836
rect 4336 16892 4400 16896
rect 4336 16836 4340 16892
rect 4340 16836 4396 16892
rect 4396 16836 4400 16892
rect 4336 16832 4400 16836
rect 4416 16892 4480 16896
rect 4416 16836 4420 16892
rect 4420 16836 4476 16892
rect 4476 16836 4480 16892
rect 4416 16832 4480 16836
rect 4496 16892 4560 16896
rect 4496 16836 4500 16892
rect 4500 16836 4556 16892
rect 4556 16836 4560 16892
rect 4496 16832 4560 16836
rect 10176 16892 10240 16896
rect 10176 16836 10180 16892
rect 10180 16836 10236 16892
rect 10236 16836 10240 16892
rect 10176 16832 10240 16836
rect 10256 16892 10320 16896
rect 10256 16836 10260 16892
rect 10260 16836 10316 16892
rect 10316 16836 10320 16892
rect 10256 16832 10320 16836
rect 10336 16892 10400 16896
rect 10336 16836 10340 16892
rect 10340 16836 10396 16892
rect 10396 16836 10400 16892
rect 10336 16832 10400 16836
rect 10416 16892 10480 16896
rect 10416 16836 10420 16892
rect 10420 16836 10476 16892
rect 10476 16836 10480 16892
rect 10416 16832 10480 16836
rect 10496 16892 10560 16896
rect 10496 16836 10500 16892
rect 10500 16836 10556 16892
rect 10556 16836 10560 16892
rect 10496 16832 10560 16836
rect 16176 16892 16240 16896
rect 16176 16836 16180 16892
rect 16180 16836 16236 16892
rect 16236 16836 16240 16892
rect 16176 16832 16240 16836
rect 16256 16892 16320 16896
rect 16256 16836 16260 16892
rect 16260 16836 16316 16892
rect 16316 16836 16320 16892
rect 16256 16832 16320 16836
rect 16336 16892 16400 16896
rect 16336 16836 16340 16892
rect 16340 16836 16396 16892
rect 16396 16836 16400 16892
rect 16336 16832 16400 16836
rect 16416 16892 16480 16896
rect 16416 16836 16420 16892
rect 16420 16836 16476 16892
rect 16476 16836 16480 16892
rect 16416 16832 16480 16836
rect 16496 16892 16560 16896
rect 16496 16836 16500 16892
rect 16500 16836 16556 16892
rect 16556 16836 16560 16892
rect 16496 16832 16560 16836
rect 22176 16892 22240 16896
rect 22176 16836 22180 16892
rect 22180 16836 22236 16892
rect 22236 16836 22240 16892
rect 22176 16832 22240 16836
rect 22256 16892 22320 16896
rect 22256 16836 22260 16892
rect 22260 16836 22316 16892
rect 22316 16836 22320 16892
rect 22256 16832 22320 16836
rect 22336 16892 22400 16896
rect 22336 16836 22340 16892
rect 22340 16836 22396 16892
rect 22396 16836 22400 16892
rect 22336 16832 22400 16836
rect 22416 16892 22480 16896
rect 22416 16836 22420 16892
rect 22420 16836 22476 16892
rect 22476 16836 22480 16892
rect 22416 16832 22480 16836
rect 22496 16892 22560 16896
rect 22496 16836 22500 16892
rect 22500 16836 22556 16892
rect 22556 16836 22560 16892
rect 22496 16832 22560 16836
rect 28176 16892 28240 16896
rect 28176 16836 28180 16892
rect 28180 16836 28236 16892
rect 28236 16836 28240 16892
rect 28176 16832 28240 16836
rect 28256 16892 28320 16896
rect 28256 16836 28260 16892
rect 28260 16836 28316 16892
rect 28316 16836 28320 16892
rect 28256 16832 28320 16836
rect 28336 16892 28400 16896
rect 28336 16836 28340 16892
rect 28340 16836 28396 16892
rect 28396 16836 28400 16892
rect 28336 16832 28400 16836
rect 28416 16892 28480 16896
rect 28416 16836 28420 16892
rect 28420 16836 28476 16892
rect 28476 16836 28480 16892
rect 28416 16832 28480 16836
rect 28496 16892 28560 16896
rect 28496 16836 28500 16892
rect 28500 16836 28556 16892
rect 28556 16836 28560 16892
rect 28496 16832 28560 16836
rect 4916 16348 4980 16352
rect 4916 16292 4920 16348
rect 4920 16292 4976 16348
rect 4976 16292 4980 16348
rect 4916 16288 4980 16292
rect 4996 16348 5060 16352
rect 4996 16292 5000 16348
rect 5000 16292 5056 16348
rect 5056 16292 5060 16348
rect 4996 16288 5060 16292
rect 5076 16348 5140 16352
rect 5076 16292 5080 16348
rect 5080 16292 5136 16348
rect 5136 16292 5140 16348
rect 5076 16288 5140 16292
rect 5156 16348 5220 16352
rect 5156 16292 5160 16348
rect 5160 16292 5216 16348
rect 5216 16292 5220 16348
rect 5156 16288 5220 16292
rect 5236 16348 5300 16352
rect 5236 16292 5240 16348
rect 5240 16292 5296 16348
rect 5296 16292 5300 16348
rect 5236 16288 5300 16292
rect 10916 16348 10980 16352
rect 10916 16292 10920 16348
rect 10920 16292 10976 16348
rect 10976 16292 10980 16348
rect 10916 16288 10980 16292
rect 10996 16348 11060 16352
rect 10996 16292 11000 16348
rect 11000 16292 11056 16348
rect 11056 16292 11060 16348
rect 10996 16288 11060 16292
rect 11076 16348 11140 16352
rect 11076 16292 11080 16348
rect 11080 16292 11136 16348
rect 11136 16292 11140 16348
rect 11076 16288 11140 16292
rect 11156 16348 11220 16352
rect 11156 16292 11160 16348
rect 11160 16292 11216 16348
rect 11216 16292 11220 16348
rect 11156 16288 11220 16292
rect 11236 16348 11300 16352
rect 11236 16292 11240 16348
rect 11240 16292 11296 16348
rect 11296 16292 11300 16348
rect 11236 16288 11300 16292
rect 16916 16348 16980 16352
rect 16916 16292 16920 16348
rect 16920 16292 16976 16348
rect 16976 16292 16980 16348
rect 16916 16288 16980 16292
rect 16996 16348 17060 16352
rect 16996 16292 17000 16348
rect 17000 16292 17056 16348
rect 17056 16292 17060 16348
rect 16996 16288 17060 16292
rect 17076 16348 17140 16352
rect 17076 16292 17080 16348
rect 17080 16292 17136 16348
rect 17136 16292 17140 16348
rect 17076 16288 17140 16292
rect 17156 16348 17220 16352
rect 17156 16292 17160 16348
rect 17160 16292 17216 16348
rect 17216 16292 17220 16348
rect 17156 16288 17220 16292
rect 17236 16348 17300 16352
rect 17236 16292 17240 16348
rect 17240 16292 17296 16348
rect 17296 16292 17300 16348
rect 17236 16288 17300 16292
rect 22916 16348 22980 16352
rect 22916 16292 22920 16348
rect 22920 16292 22976 16348
rect 22976 16292 22980 16348
rect 22916 16288 22980 16292
rect 22996 16348 23060 16352
rect 22996 16292 23000 16348
rect 23000 16292 23056 16348
rect 23056 16292 23060 16348
rect 22996 16288 23060 16292
rect 23076 16348 23140 16352
rect 23076 16292 23080 16348
rect 23080 16292 23136 16348
rect 23136 16292 23140 16348
rect 23076 16288 23140 16292
rect 23156 16348 23220 16352
rect 23156 16292 23160 16348
rect 23160 16292 23216 16348
rect 23216 16292 23220 16348
rect 23156 16288 23220 16292
rect 23236 16348 23300 16352
rect 23236 16292 23240 16348
rect 23240 16292 23296 16348
rect 23296 16292 23300 16348
rect 23236 16288 23300 16292
rect 28916 16348 28980 16352
rect 28916 16292 28920 16348
rect 28920 16292 28976 16348
rect 28976 16292 28980 16348
rect 28916 16288 28980 16292
rect 28996 16348 29060 16352
rect 28996 16292 29000 16348
rect 29000 16292 29056 16348
rect 29056 16292 29060 16348
rect 28996 16288 29060 16292
rect 29076 16348 29140 16352
rect 29076 16292 29080 16348
rect 29080 16292 29136 16348
rect 29136 16292 29140 16348
rect 29076 16288 29140 16292
rect 29156 16348 29220 16352
rect 29156 16292 29160 16348
rect 29160 16292 29216 16348
rect 29216 16292 29220 16348
rect 29156 16288 29220 16292
rect 29236 16348 29300 16352
rect 29236 16292 29240 16348
rect 29240 16292 29296 16348
rect 29296 16292 29300 16348
rect 29236 16288 29300 16292
rect 4176 15804 4240 15808
rect 4176 15748 4180 15804
rect 4180 15748 4236 15804
rect 4236 15748 4240 15804
rect 4176 15744 4240 15748
rect 4256 15804 4320 15808
rect 4256 15748 4260 15804
rect 4260 15748 4316 15804
rect 4316 15748 4320 15804
rect 4256 15744 4320 15748
rect 4336 15804 4400 15808
rect 4336 15748 4340 15804
rect 4340 15748 4396 15804
rect 4396 15748 4400 15804
rect 4336 15744 4400 15748
rect 4416 15804 4480 15808
rect 4416 15748 4420 15804
rect 4420 15748 4476 15804
rect 4476 15748 4480 15804
rect 4416 15744 4480 15748
rect 4496 15804 4560 15808
rect 4496 15748 4500 15804
rect 4500 15748 4556 15804
rect 4556 15748 4560 15804
rect 4496 15744 4560 15748
rect 10176 15804 10240 15808
rect 10176 15748 10180 15804
rect 10180 15748 10236 15804
rect 10236 15748 10240 15804
rect 10176 15744 10240 15748
rect 10256 15804 10320 15808
rect 10256 15748 10260 15804
rect 10260 15748 10316 15804
rect 10316 15748 10320 15804
rect 10256 15744 10320 15748
rect 10336 15804 10400 15808
rect 10336 15748 10340 15804
rect 10340 15748 10396 15804
rect 10396 15748 10400 15804
rect 10336 15744 10400 15748
rect 10416 15804 10480 15808
rect 10416 15748 10420 15804
rect 10420 15748 10476 15804
rect 10476 15748 10480 15804
rect 10416 15744 10480 15748
rect 10496 15804 10560 15808
rect 10496 15748 10500 15804
rect 10500 15748 10556 15804
rect 10556 15748 10560 15804
rect 10496 15744 10560 15748
rect 16176 15804 16240 15808
rect 16176 15748 16180 15804
rect 16180 15748 16236 15804
rect 16236 15748 16240 15804
rect 16176 15744 16240 15748
rect 16256 15804 16320 15808
rect 16256 15748 16260 15804
rect 16260 15748 16316 15804
rect 16316 15748 16320 15804
rect 16256 15744 16320 15748
rect 16336 15804 16400 15808
rect 16336 15748 16340 15804
rect 16340 15748 16396 15804
rect 16396 15748 16400 15804
rect 16336 15744 16400 15748
rect 16416 15804 16480 15808
rect 16416 15748 16420 15804
rect 16420 15748 16476 15804
rect 16476 15748 16480 15804
rect 16416 15744 16480 15748
rect 16496 15804 16560 15808
rect 16496 15748 16500 15804
rect 16500 15748 16556 15804
rect 16556 15748 16560 15804
rect 16496 15744 16560 15748
rect 22176 15804 22240 15808
rect 22176 15748 22180 15804
rect 22180 15748 22236 15804
rect 22236 15748 22240 15804
rect 22176 15744 22240 15748
rect 22256 15804 22320 15808
rect 22256 15748 22260 15804
rect 22260 15748 22316 15804
rect 22316 15748 22320 15804
rect 22256 15744 22320 15748
rect 22336 15804 22400 15808
rect 22336 15748 22340 15804
rect 22340 15748 22396 15804
rect 22396 15748 22400 15804
rect 22336 15744 22400 15748
rect 22416 15804 22480 15808
rect 22416 15748 22420 15804
rect 22420 15748 22476 15804
rect 22476 15748 22480 15804
rect 22416 15744 22480 15748
rect 22496 15804 22560 15808
rect 22496 15748 22500 15804
rect 22500 15748 22556 15804
rect 22556 15748 22560 15804
rect 22496 15744 22560 15748
rect 28176 15804 28240 15808
rect 28176 15748 28180 15804
rect 28180 15748 28236 15804
rect 28236 15748 28240 15804
rect 28176 15744 28240 15748
rect 28256 15804 28320 15808
rect 28256 15748 28260 15804
rect 28260 15748 28316 15804
rect 28316 15748 28320 15804
rect 28256 15744 28320 15748
rect 28336 15804 28400 15808
rect 28336 15748 28340 15804
rect 28340 15748 28396 15804
rect 28396 15748 28400 15804
rect 28336 15744 28400 15748
rect 28416 15804 28480 15808
rect 28416 15748 28420 15804
rect 28420 15748 28476 15804
rect 28476 15748 28480 15804
rect 28416 15744 28480 15748
rect 28496 15804 28560 15808
rect 28496 15748 28500 15804
rect 28500 15748 28556 15804
rect 28556 15748 28560 15804
rect 28496 15744 28560 15748
rect 4916 15260 4980 15264
rect 4916 15204 4920 15260
rect 4920 15204 4976 15260
rect 4976 15204 4980 15260
rect 4916 15200 4980 15204
rect 4996 15260 5060 15264
rect 4996 15204 5000 15260
rect 5000 15204 5056 15260
rect 5056 15204 5060 15260
rect 4996 15200 5060 15204
rect 5076 15260 5140 15264
rect 5076 15204 5080 15260
rect 5080 15204 5136 15260
rect 5136 15204 5140 15260
rect 5076 15200 5140 15204
rect 5156 15260 5220 15264
rect 5156 15204 5160 15260
rect 5160 15204 5216 15260
rect 5216 15204 5220 15260
rect 5156 15200 5220 15204
rect 5236 15260 5300 15264
rect 5236 15204 5240 15260
rect 5240 15204 5296 15260
rect 5296 15204 5300 15260
rect 5236 15200 5300 15204
rect 10916 15260 10980 15264
rect 10916 15204 10920 15260
rect 10920 15204 10976 15260
rect 10976 15204 10980 15260
rect 10916 15200 10980 15204
rect 10996 15260 11060 15264
rect 10996 15204 11000 15260
rect 11000 15204 11056 15260
rect 11056 15204 11060 15260
rect 10996 15200 11060 15204
rect 11076 15260 11140 15264
rect 11076 15204 11080 15260
rect 11080 15204 11136 15260
rect 11136 15204 11140 15260
rect 11076 15200 11140 15204
rect 11156 15260 11220 15264
rect 11156 15204 11160 15260
rect 11160 15204 11216 15260
rect 11216 15204 11220 15260
rect 11156 15200 11220 15204
rect 11236 15260 11300 15264
rect 11236 15204 11240 15260
rect 11240 15204 11296 15260
rect 11296 15204 11300 15260
rect 11236 15200 11300 15204
rect 16916 15260 16980 15264
rect 16916 15204 16920 15260
rect 16920 15204 16976 15260
rect 16976 15204 16980 15260
rect 16916 15200 16980 15204
rect 16996 15260 17060 15264
rect 16996 15204 17000 15260
rect 17000 15204 17056 15260
rect 17056 15204 17060 15260
rect 16996 15200 17060 15204
rect 17076 15260 17140 15264
rect 17076 15204 17080 15260
rect 17080 15204 17136 15260
rect 17136 15204 17140 15260
rect 17076 15200 17140 15204
rect 17156 15260 17220 15264
rect 17156 15204 17160 15260
rect 17160 15204 17216 15260
rect 17216 15204 17220 15260
rect 17156 15200 17220 15204
rect 17236 15260 17300 15264
rect 17236 15204 17240 15260
rect 17240 15204 17296 15260
rect 17296 15204 17300 15260
rect 17236 15200 17300 15204
rect 22916 15260 22980 15264
rect 22916 15204 22920 15260
rect 22920 15204 22976 15260
rect 22976 15204 22980 15260
rect 22916 15200 22980 15204
rect 22996 15260 23060 15264
rect 22996 15204 23000 15260
rect 23000 15204 23056 15260
rect 23056 15204 23060 15260
rect 22996 15200 23060 15204
rect 23076 15260 23140 15264
rect 23076 15204 23080 15260
rect 23080 15204 23136 15260
rect 23136 15204 23140 15260
rect 23076 15200 23140 15204
rect 23156 15260 23220 15264
rect 23156 15204 23160 15260
rect 23160 15204 23216 15260
rect 23216 15204 23220 15260
rect 23156 15200 23220 15204
rect 23236 15260 23300 15264
rect 23236 15204 23240 15260
rect 23240 15204 23296 15260
rect 23296 15204 23300 15260
rect 23236 15200 23300 15204
rect 28916 15260 28980 15264
rect 28916 15204 28920 15260
rect 28920 15204 28976 15260
rect 28976 15204 28980 15260
rect 28916 15200 28980 15204
rect 28996 15260 29060 15264
rect 28996 15204 29000 15260
rect 29000 15204 29056 15260
rect 29056 15204 29060 15260
rect 28996 15200 29060 15204
rect 29076 15260 29140 15264
rect 29076 15204 29080 15260
rect 29080 15204 29136 15260
rect 29136 15204 29140 15260
rect 29076 15200 29140 15204
rect 29156 15260 29220 15264
rect 29156 15204 29160 15260
rect 29160 15204 29216 15260
rect 29216 15204 29220 15260
rect 29156 15200 29220 15204
rect 29236 15260 29300 15264
rect 29236 15204 29240 15260
rect 29240 15204 29296 15260
rect 29296 15204 29300 15260
rect 29236 15200 29300 15204
rect 4176 14716 4240 14720
rect 4176 14660 4180 14716
rect 4180 14660 4236 14716
rect 4236 14660 4240 14716
rect 4176 14656 4240 14660
rect 4256 14716 4320 14720
rect 4256 14660 4260 14716
rect 4260 14660 4316 14716
rect 4316 14660 4320 14716
rect 4256 14656 4320 14660
rect 4336 14716 4400 14720
rect 4336 14660 4340 14716
rect 4340 14660 4396 14716
rect 4396 14660 4400 14716
rect 4336 14656 4400 14660
rect 4416 14716 4480 14720
rect 4416 14660 4420 14716
rect 4420 14660 4476 14716
rect 4476 14660 4480 14716
rect 4416 14656 4480 14660
rect 4496 14716 4560 14720
rect 4496 14660 4500 14716
rect 4500 14660 4556 14716
rect 4556 14660 4560 14716
rect 4496 14656 4560 14660
rect 10176 14716 10240 14720
rect 10176 14660 10180 14716
rect 10180 14660 10236 14716
rect 10236 14660 10240 14716
rect 10176 14656 10240 14660
rect 10256 14716 10320 14720
rect 10256 14660 10260 14716
rect 10260 14660 10316 14716
rect 10316 14660 10320 14716
rect 10256 14656 10320 14660
rect 10336 14716 10400 14720
rect 10336 14660 10340 14716
rect 10340 14660 10396 14716
rect 10396 14660 10400 14716
rect 10336 14656 10400 14660
rect 10416 14716 10480 14720
rect 10416 14660 10420 14716
rect 10420 14660 10476 14716
rect 10476 14660 10480 14716
rect 10416 14656 10480 14660
rect 10496 14716 10560 14720
rect 10496 14660 10500 14716
rect 10500 14660 10556 14716
rect 10556 14660 10560 14716
rect 10496 14656 10560 14660
rect 16176 14716 16240 14720
rect 16176 14660 16180 14716
rect 16180 14660 16236 14716
rect 16236 14660 16240 14716
rect 16176 14656 16240 14660
rect 16256 14716 16320 14720
rect 16256 14660 16260 14716
rect 16260 14660 16316 14716
rect 16316 14660 16320 14716
rect 16256 14656 16320 14660
rect 16336 14716 16400 14720
rect 16336 14660 16340 14716
rect 16340 14660 16396 14716
rect 16396 14660 16400 14716
rect 16336 14656 16400 14660
rect 16416 14716 16480 14720
rect 16416 14660 16420 14716
rect 16420 14660 16476 14716
rect 16476 14660 16480 14716
rect 16416 14656 16480 14660
rect 16496 14716 16560 14720
rect 16496 14660 16500 14716
rect 16500 14660 16556 14716
rect 16556 14660 16560 14716
rect 16496 14656 16560 14660
rect 22176 14716 22240 14720
rect 22176 14660 22180 14716
rect 22180 14660 22236 14716
rect 22236 14660 22240 14716
rect 22176 14656 22240 14660
rect 22256 14716 22320 14720
rect 22256 14660 22260 14716
rect 22260 14660 22316 14716
rect 22316 14660 22320 14716
rect 22256 14656 22320 14660
rect 22336 14716 22400 14720
rect 22336 14660 22340 14716
rect 22340 14660 22396 14716
rect 22396 14660 22400 14716
rect 22336 14656 22400 14660
rect 22416 14716 22480 14720
rect 22416 14660 22420 14716
rect 22420 14660 22476 14716
rect 22476 14660 22480 14716
rect 22416 14656 22480 14660
rect 22496 14716 22560 14720
rect 22496 14660 22500 14716
rect 22500 14660 22556 14716
rect 22556 14660 22560 14716
rect 22496 14656 22560 14660
rect 28176 14716 28240 14720
rect 28176 14660 28180 14716
rect 28180 14660 28236 14716
rect 28236 14660 28240 14716
rect 28176 14656 28240 14660
rect 28256 14716 28320 14720
rect 28256 14660 28260 14716
rect 28260 14660 28316 14716
rect 28316 14660 28320 14716
rect 28256 14656 28320 14660
rect 28336 14716 28400 14720
rect 28336 14660 28340 14716
rect 28340 14660 28396 14716
rect 28396 14660 28400 14716
rect 28336 14656 28400 14660
rect 28416 14716 28480 14720
rect 28416 14660 28420 14716
rect 28420 14660 28476 14716
rect 28476 14660 28480 14716
rect 28416 14656 28480 14660
rect 28496 14716 28560 14720
rect 28496 14660 28500 14716
rect 28500 14660 28556 14716
rect 28556 14660 28560 14716
rect 28496 14656 28560 14660
rect 4916 14172 4980 14176
rect 4916 14116 4920 14172
rect 4920 14116 4976 14172
rect 4976 14116 4980 14172
rect 4916 14112 4980 14116
rect 4996 14172 5060 14176
rect 4996 14116 5000 14172
rect 5000 14116 5056 14172
rect 5056 14116 5060 14172
rect 4996 14112 5060 14116
rect 5076 14172 5140 14176
rect 5076 14116 5080 14172
rect 5080 14116 5136 14172
rect 5136 14116 5140 14172
rect 5076 14112 5140 14116
rect 5156 14172 5220 14176
rect 5156 14116 5160 14172
rect 5160 14116 5216 14172
rect 5216 14116 5220 14172
rect 5156 14112 5220 14116
rect 5236 14172 5300 14176
rect 5236 14116 5240 14172
rect 5240 14116 5296 14172
rect 5296 14116 5300 14172
rect 5236 14112 5300 14116
rect 10916 14172 10980 14176
rect 10916 14116 10920 14172
rect 10920 14116 10976 14172
rect 10976 14116 10980 14172
rect 10916 14112 10980 14116
rect 10996 14172 11060 14176
rect 10996 14116 11000 14172
rect 11000 14116 11056 14172
rect 11056 14116 11060 14172
rect 10996 14112 11060 14116
rect 11076 14172 11140 14176
rect 11076 14116 11080 14172
rect 11080 14116 11136 14172
rect 11136 14116 11140 14172
rect 11076 14112 11140 14116
rect 11156 14172 11220 14176
rect 11156 14116 11160 14172
rect 11160 14116 11216 14172
rect 11216 14116 11220 14172
rect 11156 14112 11220 14116
rect 11236 14172 11300 14176
rect 11236 14116 11240 14172
rect 11240 14116 11296 14172
rect 11296 14116 11300 14172
rect 11236 14112 11300 14116
rect 16916 14172 16980 14176
rect 16916 14116 16920 14172
rect 16920 14116 16976 14172
rect 16976 14116 16980 14172
rect 16916 14112 16980 14116
rect 16996 14172 17060 14176
rect 16996 14116 17000 14172
rect 17000 14116 17056 14172
rect 17056 14116 17060 14172
rect 16996 14112 17060 14116
rect 17076 14172 17140 14176
rect 17076 14116 17080 14172
rect 17080 14116 17136 14172
rect 17136 14116 17140 14172
rect 17076 14112 17140 14116
rect 17156 14172 17220 14176
rect 17156 14116 17160 14172
rect 17160 14116 17216 14172
rect 17216 14116 17220 14172
rect 17156 14112 17220 14116
rect 17236 14172 17300 14176
rect 17236 14116 17240 14172
rect 17240 14116 17296 14172
rect 17296 14116 17300 14172
rect 17236 14112 17300 14116
rect 22916 14172 22980 14176
rect 22916 14116 22920 14172
rect 22920 14116 22976 14172
rect 22976 14116 22980 14172
rect 22916 14112 22980 14116
rect 22996 14172 23060 14176
rect 22996 14116 23000 14172
rect 23000 14116 23056 14172
rect 23056 14116 23060 14172
rect 22996 14112 23060 14116
rect 23076 14172 23140 14176
rect 23076 14116 23080 14172
rect 23080 14116 23136 14172
rect 23136 14116 23140 14172
rect 23076 14112 23140 14116
rect 23156 14172 23220 14176
rect 23156 14116 23160 14172
rect 23160 14116 23216 14172
rect 23216 14116 23220 14172
rect 23156 14112 23220 14116
rect 23236 14172 23300 14176
rect 23236 14116 23240 14172
rect 23240 14116 23296 14172
rect 23296 14116 23300 14172
rect 23236 14112 23300 14116
rect 28916 14172 28980 14176
rect 28916 14116 28920 14172
rect 28920 14116 28976 14172
rect 28976 14116 28980 14172
rect 28916 14112 28980 14116
rect 28996 14172 29060 14176
rect 28996 14116 29000 14172
rect 29000 14116 29056 14172
rect 29056 14116 29060 14172
rect 28996 14112 29060 14116
rect 29076 14172 29140 14176
rect 29076 14116 29080 14172
rect 29080 14116 29136 14172
rect 29136 14116 29140 14172
rect 29076 14112 29140 14116
rect 29156 14172 29220 14176
rect 29156 14116 29160 14172
rect 29160 14116 29216 14172
rect 29216 14116 29220 14172
rect 29156 14112 29220 14116
rect 29236 14172 29300 14176
rect 29236 14116 29240 14172
rect 29240 14116 29296 14172
rect 29296 14116 29300 14172
rect 29236 14112 29300 14116
rect 4176 13628 4240 13632
rect 4176 13572 4180 13628
rect 4180 13572 4236 13628
rect 4236 13572 4240 13628
rect 4176 13568 4240 13572
rect 4256 13628 4320 13632
rect 4256 13572 4260 13628
rect 4260 13572 4316 13628
rect 4316 13572 4320 13628
rect 4256 13568 4320 13572
rect 4336 13628 4400 13632
rect 4336 13572 4340 13628
rect 4340 13572 4396 13628
rect 4396 13572 4400 13628
rect 4336 13568 4400 13572
rect 4416 13628 4480 13632
rect 4416 13572 4420 13628
rect 4420 13572 4476 13628
rect 4476 13572 4480 13628
rect 4416 13568 4480 13572
rect 4496 13628 4560 13632
rect 4496 13572 4500 13628
rect 4500 13572 4556 13628
rect 4556 13572 4560 13628
rect 4496 13568 4560 13572
rect 10176 13628 10240 13632
rect 10176 13572 10180 13628
rect 10180 13572 10236 13628
rect 10236 13572 10240 13628
rect 10176 13568 10240 13572
rect 10256 13628 10320 13632
rect 10256 13572 10260 13628
rect 10260 13572 10316 13628
rect 10316 13572 10320 13628
rect 10256 13568 10320 13572
rect 10336 13628 10400 13632
rect 10336 13572 10340 13628
rect 10340 13572 10396 13628
rect 10396 13572 10400 13628
rect 10336 13568 10400 13572
rect 10416 13628 10480 13632
rect 10416 13572 10420 13628
rect 10420 13572 10476 13628
rect 10476 13572 10480 13628
rect 10416 13568 10480 13572
rect 10496 13628 10560 13632
rect 10496 13572 10500 13628
rect 10500 13572 10556 13628
rect 10556 13572 10560 13628
rect 10496 13568 10560 13572
rect 16176 13628 16240 13632
rect 16176 13572 16180 13628
rect 16180 13572 16236 13628
rect 16236 13572 16240 13628
rect 16176 13568 16240 13572
rect 16256 13628 16320 13632
rect 16256 13572 16260 13628
rect 16260 13572 16316 13628
rect 16316 13572 16320 13628
rect 16256 13568 16320 13572
rect 16336 13628 16400 13632
rect 16336 13572 16340 13628
rect 16340 13572 16396 13628
rect 16396 13572 16400 13628
rect 16336 13568 16400 13572
rect 16416 13628 16480 13632
rect 16416 13572 16420 13628
rect 16420 13572 16476 13628
rect 16476 13572 16480 13628
rect 16416 13568 16480 13572
rect 16496 13628 16560 13632
rect 16496 13572 16500 13628
rect 16500 13572 16556 13628
rect 16556 13572 16560 13628
rect 16496 13568 16560 13572
rect 22176 13628 22240 13632
rect 22176 13572 22180 13628
rect 22180 13572 22236 13628
rect 22236 13572 22240 13628
rect 22176 13568 22240 13572
rect 22256 13628 22320 13632
rect 22256 13572 22260 13628
rect 22260 13572 22316 13628
rect 22316 13572 22320 13628
rect 22256 13568 22320 13572
rect 22336 13628 22400 13632
rect 22336 13572 22340 13628
rect 22340 13572 22396 13628
rect 22396 13572 22400 13628
rect 22336 13568 22400 13572
rect 22416 13628 22480 13632
rect 22416 13572 22420 13628
rect 22420 13572 22476 13628
rect 22476 13572 22480 13628
rect 22416 13568 22480 13572
rect 22496 13628 22560 13632
rect 22496 13572 22500 13628
rect 22500 13572 22556 13628
rect 22556 13572 22560 13628
rect 22496 13568 22560 13572
rect 28176 13628 28240 13632
rect 28176 13572 28180 13628
rect 28180 13572 28236 13628
rect 28236 13572 28240 13628
rect 28176 13568 28240 13572
rect 28256 13628 28320 13632
rect 28256 13572 28260 13628
rect 28260 13572 28316 13628
rect 28316 13572 28320 13628
rect 28256 13568 28320 13572
rect 28336 13628 28400 13632
rect 28336 13572 28340 13628
rect 28340 13572 28396 13628
rect 28396 13572 28400 13628
rect 28336 13568 28400 13572
rect 28416 13628 28480 13632
rect 28416 13572 28420 13628
rect 28420 13572 28476 13628
rect 28476 13572 28480 13628
rect 28416 13568 28480 13572
rect 28496 13628 28560 13632
rect 28496 13572 28500 13628
rect 28500 13572 28556 13628
rect 28556 13572 28560 13628
rect 28496 13568 28560 13572
rect 4916 13084 4980 13088
rect 4916 13028 4920 13084
rect 4920 13028 4976 13084
rect 4976 13028 4980 13084
rect 4916 13024 4980 13028
rect 4996 13084 5060 13088
rect 4996 13028 5000 13084
rect 5000 13028 5056 13084
rect 5056 13028 5060 13084
rect 4996 13024 5060 13028
rect 5076 13084 5140 13088
rect 5076 13028 5080 13084
rect 5080 13028 5136 13084
rect 5136 13028 5140 13084
rect 5076 13024 5140 13028
rect 5156 13084 5220 13088
rect 5156 13028 5160 13084
rect 5160 13028 5216 13084
rect 5216 13028 5220 13084
rect 5156 13024 5220 13028
rect 5236 13084 5300 13088
rect 5236 13028 5240 13084
rect 5240 13028 5296 13084
rect 5296 13028 5300 13084
rect 5236 13024 5300 13028
rect 10916 13084 10980 13088
rect 10916 13028 10920 13084
rect 10920 13028 10976 13084
rect 10976 13028 10980 13084
rect 10916 13024 10980 13028
rect 10996 13084 11060 13088
rect 10996 13028 11000 13084
rect 11000 13028 11056 13084
rect 11056 13028 11060 13084
rect 10996 13024 11060 13028
rect 11076 13084 11140 13088
rect 11076 13028 11080 13084
rect 11080 13028 11136 13084
rect 11136 13028 11140 13084
rect 11076 13024 11140 13028
rect 11156 13084 11220 13088
rect 11156 13028 11160 13084
rect 11160 13028 11216 13084
rect 11216 13028 11220 13084
rect 11156 13024 11220 13028
rect 11236 13084 11300 13088
rect 11236 13028 11240 13084
rect 11240 13028 11296 13084
rect 11296 13028 11300 13084
rect 11236 13024 11300 13028
rect 16916 13084 16980 13088
rect 16916 13028 16920 13084
rect 16920 13028 16976 13084
rect 16976 13028 16980 13084
rect 16916 13024 16980 13028
rect 16996 13084 17060 13088
rect 16996 13028 17000 13084
rect 17000 13028 17056 13084
rect 17056 13028 17060 13084
rect 16996 13024 17060 13028
rect 17076 13084 17140 13088
rect 17076 13028 17080 13084
rect 17080 13028 17136 13084
rect 17136 13028 17140 13084
rect 17076 13024 17140 13028
rect 17156 13084 17220 13088
rect 17156 13028 17160 13084
rect 17160 13028 17216 13084
rect 17216 13028 17220 13084
rect 17156 13024 17220 13028
rect 17236 13084 17300 13088
rect 17236 13028 17240 13084
rect 17240 13028 17296 13084
rect 17296 13028 17300 13084
rect 17236 13024 17300 13028
rect 22916 13084 22980 13088
rect 22916 13028 22920 13084
rect 22920 13028 22976 13084
rect 22976 13028 22980 13084
rect 22916 13024 22980 13028
rect 22996 13084 23060 13088
rect 22996 13028 23000 13084
rect 23000 13028 23056 13084
rect 23056 13028 23060 13084
rect 22996 13024 23060 13028
rect 23076 13084 23140 13088
rect 23076 13028 23080 13084
rect 23080 13028 23136 13084
rect 23136 13028 23140 13084
rect 23076 13024 23140 13028
rect 23156 13084 23220 13088
rect 23156 13028 23160 13084
rect 23160 13028 23216 13084
rect 23216 13028 23220 13084
rect 23156 13024 23220 13028
rect 23236 13084 23300 13088
rect 23236 13028 23240 13084
rect 23240 13028 23296 13084
rect 23296 13028 23300 13084
rect 23236 13024 23300 13028
rect 28916 13084 28980 13088
rect 28916 13028 28920 13084
rect 28920 13028 28976 13084
rect 28976 13028 28980 13084
rect 28916 13024 28980 13028
rect 28996 13084 29060 13088
rect 28996 13028 29000 13084
rect 29000 13028 29056 13084
rect 29056 13028 29060 13084
rect 28996 13024 29060 13028
rect 29076 13084 29140 13088
rect 29076 13028 29080 13084
rect 29080 13028 29136 13084
rect 29136 13028 29140 13084
rect 29076 13024 29140 13028
rect 29156 13084 29220 13088
rect 29156 13028 29160 13084
rect 29160 13028 29216 13084
rect 29216 13028 29220 13084
rect 29156 13024 29220 13028
rect 29236 13084 29300 13088
rect 29236 13028 29240 13084
rect 29240 13028 29296 13084
rect 29296 13028 29300 13084
rect 29236 13024 29300 13028
rect 12940 12684 13004 12748
rect 19380 12684 19444 12748
rect 4176 12540 4240 12544
rect 4176 12484 4180 12540
rect 4180 12484 4236 12540
rect 4236 12484 4240 12540
rect 4176 12480 4240 12484
rect 4256 12540 4320 12544
rect 4256 12484 4260 12540
rect 4260 12484 4316 12540
rect 4316 12484 4320 12540
rect 4256 12480 4320 12484
rect 4336 12540 4400 12544
rect 4336 12484 4340 12540
rect 4340 12484 4396 12540
rect 4396 12484 4400 12540
rect 4336 12480 4400 12484
rect 4416 12540 4480 12544
rect 4416 12484 4420 12540
rect 4420 12484 4476 12540
rect 4476 12484 4480 12540
rect 4416 12480 4480 12484
rect 4496 12540 4560 12544
rect 4496 12484 4500 12540
rect 4500 12484 4556 12540
rect 4556 12484 4560 12540
rect 4496 12480 4560 12484
rect 10176 12540 10240 12544
rect 10176 12484 10180 12540
rect 10180 12484 10236 12540
rect 10236 12484 10240 12540
rect 10176 12480 10240 12484
rect 10256 12540 10320 12544
rect 10256 12484 10260 12540
rect 10260 12484 10316 12540
rect 10316 12484 10320 12540
rect 10256 12480 10320 12484
rect 10336 12540 10400 12544
rect 10336 12484 10340 12540
rect 10340 12484 10396 12540
rect 10396 12484 10400 12540
rect 10336 12480 10400 12484
rect 10416 12540 10480 12544
rect 10416 12484 10420 12540
rect 10420 12484 10476 12540
rect 10476 12484 10480 12540
rect 10416 12480 10480 12484
rect 10496 12540 10560 12544
rect 10496 12484 10500 12540
rect 10500 12484 10556 12540
rect 10556 12484 10560 12540
rect 10496 12480 10560 12484
rect 16176 12540 16240 12544
rect 16176 12484 16180 12540
rect 16180 12484 16236 12540
rect 16236 12484 16240 12540
rect 16176 12480 16240 12484
rect 16256 12540 16320 12544
rect 16256 12484 16260 12540
rect 16260 12484 16316 12540
rect 16316 12484 16320 12540
rect 16256 12480 16320 12484
rect 16336 12540 16400 12544
rect 16336 12484 16340 12540
rect 16340 12484 16396 12540
rect 16396 12484 16400 12540
rect 16336 12480 16400 12484
rect 16416 12540 16480 12544
rect 16416 12484 16420 12540
rect 16420 12484 16476 12540
rect 16476 12484 16480 12540
rect 16416 12480 16480 12484
rect 16496 12540 16560 12544
rect 16496 12484 16500 12540
rect 16500 12484 16556 12540
rect 16556 12484 16560 12540
rect 16496 12480 16560 12484
rect 22176 12540 22240 12544
rect 22176 12484 22180 12540
rect 22180 12484 22236 12540
rect 22236 12484 22240 12540
rect 22176 12480 22240 12484
rect 22256 12540 22320 12544
rect 22256 12484 22260 12540
rect 22260 12484 22316 12540
rect 22316 12484 22320 12540
rect 22256 12480 22320 12484
rect 22336 12540 22400 12544
rect 22336 12484 22340 12540
rect 22340 12484 22396 12540
rect 22396 12484 22400 12540
rect 22336 12480 22400 12484
rect 22416 12540 22480 12544
rect 22416 12484 22420 12540
rect 22420 12484 22476 12540
rect 22476 12484 22480 12540
rect 22416 12480 22480 12484
rect 22496 12540 22560 12544
rect 22496 12484 22500 12540
rect 22500 12484 22556 12540
rect 22556 12484 22560 12540
rect 22496 12480 22560 12484
rect 28176 12540 28240 12544
rect 28176 12484 28180 12540
rect 28180 12484 28236 12540
rect 28236 12484 28240 12540
rect 28176 12480 28240 12484
rect 28256 12540 28320 12544
rect 28256 12484 28260 12540
rect 28260 12484 28316 12540
rect 28316 12484 28320 12540
rect 28256 12480 28320 12484
rect 28336 12540 28400 12544
rect 28336 12484 28340 12540
rect 28340 12484 28396 12540
rect 28396 12484 28400 12540
rect 28336 12480 28400 12484
rect 28416 12540 28480 12544
rect 28416 12484 28420 12540
rect 28420 12484 28476 12540
rect 28476 12484 28480 12540
rect 28416 12480 28480 12484
rect 28496 12540 28560 12544
rect 28496 12484 28500 12540
rect 28500 12484 28556 12540
rect 28556 12484 28560 12540
rect 28496 12480 28560 12484
rect 4916 11996 4980 12000
rect 4916 11940 4920 11996
rect 4920 11940 4976 11996
rect 4976 11940 4980 11996
rect 4916 11936 4980 11940
rect 4996 11996 5060 12000
rect 4996 11940 5000 11996
rect 5000 11940 5056 11996
rect 5056 11940 5060 11996
rect 4996 11936 5060 11940
rect 5076 11996 5140 12000
rect 5076 11940 5080 11996
rect 5080 11940 5136 11996
rect 5136 11940 5140 11996
rect 5076 11936 5140 11940
rect 5156 11996 5220 12000
rect 5156 11940 5160 11996
rect 5160 11940 5216 11996
rect 5216 11940 5220 11996
rect 5156 11936 5220 11940
rect 5236 11996 5300 12000
rect 5236 11940 5240 11996
rect 5240 11940 5296 11996
rect 5296 11940 5300 11996
rect 5236 11936 5300 11940
rect 10916 11996 10980 12000
rect 10916 11940 10920 11996
rect 10920 11940 10976 11996
rect 10976 11940 10980 11996
rect 10916 11936 10980 11940
rect 10996 11996 11060 12000
rect 10996 11940 11000 11996
rect 11000 11940 11056 11996
rect 11056 11940 11060 11996
rect 10996 11936 11060 11940
rect 11076 11996 11140 12000
rect 11076 11940 11080 11996
rect 11080 11940 11136 11996
rect 11136 11940 11140 11996
rect 11076 11936 11140 11940
rect 11156 11996 11220 12000
rect 11156 11940 11160 11996
rect 11160 11940 11216 11996
rect 11216 11940 11220 11996
rect 11156 11936 11220 11940
rect 11236 11996 11300 12000
rect 11236 11940 11240 11996
rect 11240 11940 11296 11996
rect 11296 11940 11300 11996
rect 11236 11936 11300 11940
rect 16916 11996 16980 12000
rect 16916 11940 16920 11996
rect 16920 11940 16976 11996
rect 16976 11940 16980 11996
rect 16916 11936 16980 11940
rect 16996 11996 17060 12000
rect 16996 11940 17000 11996
rect 17000 11940 17056 11996
rect 17056 11940 17060 11996
rect 16996 11936 17060 11940
rect 17076 11996 17140 12000
rect 17076 11940 17080 11996
rect 17080 11940 17136 11996
rect 17136 11940 17140 11996
rect 17076 11936 17140 11940
rect 17156 11996 17220 12000
rect 17156 11940 17160 11996
rect 17160 11940 17216 11996
rect 17216 11940 17220 11996
rect 17156 11936 17220 11940
rect 17236 11996 17300 12000
rect 17236 11940 17240 11996
rect 17240 11940 17296 11996
rect 17296 11940 17300 11996
rect 17236 11936 17300 11940
rect 22916 11996 22980 12000
rect 22916 11940 22920 11996
rect 22920 11940 22976 11996
rect 22976 11940 22980 11996
rect 22916 11936 22980 11940
rect 22996 11996 23060 12000
rect 22996 11940 23000 11996
rect 23000 11940 23056 11996
rect 23056 11940 23060 11996
rect 22996 11936 23060 11940
rect 23076 11996 23140 12000
rect 23076 11940 23080 11996
rect 23080 11940 23136 11996
rect 23136 11940 23140 11996
rect 23076 11936 23140 11940
rect 23156 11996 23220 12000
rect 23156 11940 23160 11996
rect 23160 11940 23216 11996
rect 23216 11940 23220 11996
rect 23156 11936 23220 11940
rect 23236 11996 23300 12000
rect 23236 11940 23240 11996
rect 23240 11940 23296 11996
rect 23296 11940 23300 11996
rect 23236 11936 23300 11940
rect 28916 11996 28980 12000
rect 28916 11940 28920 11996
rect 28920 11940 28976 11996
rect 28976 11940 28980 11996
rect 28916 11936 28980 11940
rect 28996 11996 29060 12000
rect 28996 11940 29000 11996
rect 29000 11940 29056 11996
rect 29056 11940 29060 11996
rect 28996 11936 29060 11940
rect 29076 11996 29140 12000
rect 29076 11940 29080 11996
rect 29080 11940 29136 11996
rect 29136 11940 29140 11996
rect 29076 11936 29140 11940
rect 29156 11996 29220 12000
rect 29156 11940 29160 11996
rect 29160 11940 29216 11996
rect 29216 11940 29220 11996
rect 29156 11936 29220 11940
rect 29236 11996 29300 12000
rect 29236 11940 29240 11996
rect 29240 11940 29296 11996
rect 29296 11940 29300 11996
rect 29236 11936 29300 11940
rect 4176 11452 4240 11456
rect 4176 11396 4180 11452
rect 4180 11396 4236 11452
rect 4236 11396 4240 11452
rect 4176 11392 4240 11396
rect 4256 11452 4320 11456
rect 4256 11396 4260 11452
rect 4260 11396 4316 11452
rect 4316 11396 4320 11452
rect 4256 11392 4320 11396
rect 4336 11452 4400 11456
rect 4336 11396 4340 11452
rect 4340 11396 4396 11452
rect 4396 11396 4400 11452
rect 4336 11392 4400 11396
rect 4416 11452 4480 11456
rect 4416 11396 4420 11452
rect 4420 11396 4476 11452
rect 4476 11396 4480 11452
rect 4416 11392 4480 11396
rect 4496 11452 4560 11456
rect 4496 11396 4500 11452
rect 4500 11396 4556 11452
rect 4556 11396 4560 11452
rect 4496 11392 4560 11396
rect 10176 11452 10240 11456
rect 10176 11396 10180 11452
rect 10180 11396 10236 11452
rect 10236 11396 10240 11452
rect 10176 11392 10240 11396
rect 10256 11452 10320 11456
rect 10256 11396 10260 11452
rect 10260 11396 10316 11452
rect 10316 11396 10320 11452
rect 10256 11392 10320 11396
rect 10336 11452 10400 11456
rect 10336 11396 10340 11452
rect 10340 11396 10396 11452
rect 10396 11396 10400 11452
rect 10336 11392 10400 11396
rect 10416 11452 10480 11456
rect 10416 11396 10420 11452
rect 10420 11396 10476 11452
rect 10476 11396 10480 11452
rect 10416 11392 10480 11396
rect 10496 11452 10560 11456
rect 10496 11396 10500 11452
rect 10500 11396 10556 11452
rect 10556 11396 10560 11452
rect 10496 11392 10560 11396
rect 16176 11452 16240 11456
rect 16176 11396 16180 11452
rect 16180 11396 16236 11452
rect 16236 11396 16240 11452
rect 16176 11392 16240 11396
rect 16256 11452 16320 11456
rect 16256 11396 16260 11452
rect 16260 11396 16316 11452
rect 16316 11396 16320 11452
rect 16256 11392 16320 11396
rect 16336 11452 16400 11456
rect 16336 11396 16340 11452
rect 16340 11396 16396 11452
rect 16396 11396 16400 11452
rect 16336 11392 16400 11396
rect 16416 11452 16480 11456
rect 16416 11396 16420 11452
rect 16420 11396 16476 11452
rect 16476 11396 16480 11452
rect 16416 11392 16480 11396
rect 16496 11452 16560 11456
rect 16496 11396 16500 11452
rect 16500 11396 16556 11452
rect 16556 11396 16560 11452
rect 16496 11392 16560 11396
rect 22176 11452 22240 11456
rect 22176 11396 22180 11452
rect 22180 11396 22236 11452
rect 22236 11396 22240 11452
rect 22176 11392 22240 11396
rect 22256 11452 22320 11456
rect 22256 11396 22260 11452
rect 22260 11396 22316 11452
rect 22316 11396 22320 11452
rect 22256 11392 22320 11396
rect 22336 11452 22400 11456
rect 22336 11396 22340 11452
rect 22340 11396 22396 11452
rect 22396 11396 22400 11452
rect 22336 11392 22400 11396
rect 22416 11452 22480 11456
rect 22416 11396 22420 11452
rect 22420 11396 22476 11452
rect 22476 11396 22480 11452
rect 22416 11392 22480 11396
rect 22496 11452 22560 11456
rect 22496 11396 22500 11452
rect 22500 11396 22556 11452
rect 22556 11396 22560 11452
rect 22496 11392 22560 11396
rect 28176 11452 28240 11456
rect 28176 11396 28180 11452
rect 28180 11396 28236 11452
rect 28236 11396 28240 11452
rect 28176 11392 28240 11396
rect 28256 11452 28320 11456
rect 28256 11396 28260 11452
rect 28260 11396 28316 11452
rect 28316 11396 28320 11452
rect 28256 11392 28320 11396
rect 28336 11452 28400 11456
rect 28336 11396 28340 11452
rect 28340 11396 28396 11452
rect 28396 11396 28400 11452
rect 28336 11392 28400 11396
rect 28416 11452 28480 11456
rect 28416 11396 28420 11452
rect 28420 11396 28476 11452
rect 28476 11396 28480 11452
rect 28416 11392 28480 11396
rect 28496 11452 28560 11456
rect 28496 11396 28500 11452
rect 28500 11396 28556 11452
rect 28556 11396 28560 11452
rect 28496 11392 28560 11396
rect 12940 11384 13004 11388
rect 12940 11328 12990 11384
rect 12990 11328 13004 11384
rect 12940 11324 13004 11328
rect 4916 10908 4980 10912
rect 4916 10852 4920 10908
rect 4920 10852 4976 10908
rect 4976 10852 4980 10908
rect 4916 10848 4980 10852
rect 4996 10908 5060 10912
rect 4996 10852 5000 10908
rect 5000 10852 5056 10908
rect 5056 10852 5060 10908
rect 4996 10848 5060 10852
rect 5076 10908 5140 10912
rect 5076 10852 5080 10908
rect 5080 10852 5136 10908
rect 5136 10852 5140 10908
rect 5076 10848 5140 10852
rect 5156 10908 5220 10912
rect 5156 10852 5160 10908
rect 5160 10852 5216 10908
rect 5216 10852 5220 10908
rect 5156 10848 5220 10852
rect 5236 10908 5300 10912
rect 5236 10852 5240 10908
rect 5240 10852 5296 10908
rect 5296 10852 5300 10908
rect 5236 10848 5300 10852
rect 10916 10908 10980 10912
rect 10916 10852 10920 10908
rect 10920 10852 10976 10908
rect 10976 10852 10980 10908
rect 10916 10848 10980 10852
rect 10996 10908 11060 10912
rect 10996 10852 11000 10908
rect 11000 10852 11056 10908
rect 11056 10852 11060 10908
rect 10996 10848 11060 10852
rect 11076 10908 11140 10912
rect 11076 10852 11080 10908
rect 11080 10852 11136 10908
rect 11136 10852 11140 10908
rect 11076 10848 11140 10852
rect 11156 10908 11220 10912
rect 11156 10852 11160 10908
rect 11160 10852 11216 10908
rect 11216 10852 11220 10908
rect 11156 10848 11220 10852
rect 11236 10908 11300 10912
rect 11236 10852 11240 10908
rect 11240 10852 11296 10908
rect 11296 10852 11300 10908
rect 11236 10848 11300 10852
rect 16916 10908 16980 10912
rect 16916 10852 16920 10908
rect 16920 10852 16976 10908
rect 16976 10852 16980 10908
rect 16916 10848 16980 10852
rect 16996 10908 17060 10912
rect 16996 10852 17000 10908
rect 17000 10852 17056 10908
rect 17056 10852 17060 10908
rect 16996 10848 17060 10852
rect 17076 10908 17140 10912
rect 17076 10852 17080 10908
rect 17080 10852 17136 10908
rect 17136 10852 17140 10908
rect 17076 10848 17140 10852
rect 17156 10908 17220 10912
rect 17156 10852 17160 10908
rect 17160 10852 17216 10908
rect 17216 10852 17220 10908
rect 17156 10848 17220 10852
rect 17236 10908 17300 10912
rect 17236 10852 17240 10908
rect 17240 10852 17296 10908
rect 17296 10852 17300 10908
rect 17236 10848 17300 10852
rect 22916 10908 22980 10912
rect 22916 10852 22920 10908
rect 22920 10852 22976 10908
rect 22976 10852 22980 10908
rect 22916 10848 22980 10852
rect 22996 10908 23060 10912
rect 22996 10852 23000 10908
rect 23000 10852 23056 10908
rect 23056 10852 23060 10908
rect 22996 10848 23060 10852
rect 23076 10908 23140 10912
rect 23076 10852 23080 10908
rect 23080 10852 23136 10908
rect 23136 10852 23140 10908
rect 23076 10848 23140 10852
rect 23156 10908 23220 10912
rect 23156 10852 23160 10908
rect 23160 10852 23216 10908
rect 23216 10852 23220 10908
rect 23156 10848 23220 10852
rect 23236 10908 23300 10912
rect 23236 10852 23240 10908
rect 23240 10852 23296 10908
rect 23296 10852 23300 10908
rect 23236 10848 23300 10852
rect 28916 10908 28980 10912
rect 28916 10852 28920 10908
rect 28920 10852 28976 10908
rect 28976 10852 28980 10908
rect 28916 10848 28980 10852
rect 28996 10908 29060 10912
rect 28996 10852 29000 10908
rect 29000 10852 29056 10908
rect 29056 10852 29060 10908
rect 28996 10848 29060 10852
rect 29076 10908 29140 10912
rect 29076 10852 29080 10908
rect 29080 10852 29136 10908
rect 29136 10852 29140 10908
rect 29076 10848 29140 10852
rect 29156 10908 29220 10912
rect 29156 10852 29160 10908
rect 29160 10852 29216 10908
rect 29216 10852 29220 10908
rect 29156 10848 29220 10852
rect 29236 10908 29300 10912
rect 29236 10852 29240 10908
rect 29240 10852 29296 10908
rect 29296 10852 29300 10908
rect 29236 10848 29300 10852
rect 4176 10364 4240 10368
rect 4176 10308 4180 10364
rect 4180 10308 4236 10364
rect 4236 10308 4240 10364
rect 4176 10304 4240 10308
rect 4256 10364 4320 10368
rect 4256 10308 4260 10364
rect 4260 10308 4316 10364
rect 4316 10308 4320 10364
rect 4256 10304 4320 10308
rect 4336 10364 4400 10368
rect 4336 10308 4340 10364
rect 4340 10308 4396 10364
rect 4396 10308 4400 10364
rect 4336 10304 4400 10308
rect 4416 10364 4480 10368
rect 4416 10308 4420 10364
rect 4420 10308 4476 10364
rect 4476 10308 4480 10364
rect 4416 10304 4480 10308
rect 4496 10364 4560 10368
rect 4496 10308 4500 10364
rect 4500 10308 4556 10364
rect 4556 10308 4560 10364
rect 4496 10304 4560 10308
rect 10176 10364 10240 10368
rect 10176 10308 10180 10364
rect 10180 10308 10236 10364
rect 10236 10308 10240 10364
rect 10176 10304 10240 10308
rect 10256 10364 10320 10368
rect 10256 10308 10260 10364
rect 10260 10308 10316 10364
rect 10316 10308 10320 10364
rect 10256 10304 10320 10308
rect 10336 10364 10400 10368
rect 10336 10308 10340 10364
rect 10340 10308 10396 10364
rect 10396 10308 10400 10364
rect 10336 10304 10400 10308
rect 10416 10364 10480 10368
rect 10416 10308 10420 10364
rect 10420 10308 10476 10364
rect 10476 10308 10480 10364
rect 10416 10304 10480 10308
rect 10496 10364 10560 10368
rect 10496 10308 10500 10364
rect 10500 10308 10556 10364
rect 10556 10308 10560 10364
rect 10496 10304 10560 10308
rect 16176 10364 16240 10368
rect 16176 10308 16180 10364
rect 16180 10308 16236 10364
rect 16236 10308 16240 10364
rect 16176 10304 16240 10308
rect 16256 10364 16320 10368
rect 16256 10308 16260 10364
rect 16260 10308 16316 10364
rect 16316 10308 16320 10364
rect 16256 10304 16320 10308
rect 16336 10364 16400 10368
rect 16336 10308 16340 10364
rect 16340 10308 16396 10364
rect 16396 10308 16400 10364
rect 16336 10304 16400 10308
rect 16416 10364 16480 10368
rect 16416 10308 16420 10364
rect 16420 10308 16476 10364
rect 16476 10308 16480 10364
rect 16416 10304 16480 10308
rect 16496 10364 16560 10368
rect 16496 10308 16500 10364
rect 16500 10308 16556 10364
rect 16556 10308 16560 10364
rect 16496 10304 16560 10308
rect 22176 10364 22240 10368
rect 22176 10308 22180 10364
rect 22180 10308 22236 10364
rect 22236 10308 22240 10364
rect 22176 10304 22240 10308
rect 22256 10364 22320 10368
rect 22256 10308 22260 10364
rect 22260 10308 22316 10364
rect 22316 10308 22320 10364
rect 22256 10304 22320 10308
rect 22336 10364 22400 10368
rect 22336 10308 22340 10364
rect 22340 10308 22396 10364
rect 22396 10308 22400 10364
rect 22336 10304 22400 10308
rect 22416 10364 22480 10368
rect 22416 10308 22420 10364
rect 22420 10308 22476 10364
rect 22476 10308 22480 10364
rect 22416 10304 22480 10308
rect 22496 10364 22560 10368
rect 22496 10308 22500 10364
rect 22500 10308 22556 10364
rect 22556 10308 22560 10364
rect 22496 10304 22560 10308
rect 28176 10364 28240 10368
rect 28176 10308 28180 10364
rect 28180 10308 28236 10364
rect 28236 10308 28240 10364
rect 28176 10304 28240 10308
rect 28256 10364 28320 10368
rect 28256 10308 28260 10364
rect 28260 10308 28316 10364
rect 28316 10308 28320 10364
rect 28256 10304 28320 10308
rect 28336 10364 28400 10368
rect 28336 10308 28340 10364
rect 28340 10308 28396 10364
rect 28396 10308 28400 10364
rect 28336 10304 28400 10308
rect 28416 10364 28480 10368
rect 28416 10308 28420 10364
rect 28420 10308 28476 10364
rect 28476 10308 28480 10364
rect 28416 10304 28480 10308
rect 28496 10364 28560 10368
rect 28496 10308 28500 10364
rect 28500 10308 28556 10364
rect 28556 10308 28560 10364
rect 28496 10304 28560 10308
rect 4916 9820 4980 9824
rect 4916 9764 4920 9820
rect 4920 9764 4976 9820
rect 4976 9764 4980 9820
rect 4916 9760 4980 9764
rect 4996 9820 5060 9824
rect 4996 9764 5000 9820
rect 5000 9764 5056 9820
rect 5056 9764 5060 9820
rect 4996 9760 5060 9764
rect 5076 9820 5140 9824
rect 5076 9764 5080 9820
rect 5080 9764 5136 9820
rect 5136 9764 5140 9820
rect 5076 9760 5140 9764
rect 5156 9820 5220 9824
rect 5156 9764 5160 9820
rect 5160 9764 5216 9820
rect 5216 9764 5220 9820
rect 5156 9760 5220 9764
rect 5236 9820 5300 9824
rect 5236 9764 5240 9820
rect 5240 9764 5296 9820
rect 5296 9764 5300 9820
rect 5236 9760 5300 9764
rect 10916 9820 10980 9824
rect 10916 9764 10920 9820
rect 10920 9764 10976 9820
rect 10976 9764 10980 9820
rect 10916 9760 10980 9764
rect 10996 9820 11060 9824
rect 10996 9764 11000 9820
rect 11000 9764 11056 9820
rect 11056 9764 11060 9820
rect 10996 9760 11060 9764
rect 11076 9820 11140 9824
rect 11076 9764 11080 9820
rect 11080 9764 11136 9820
rect 11136 9764 11140 9820
rect 11076 9760 11140 9764
rect 11156 9820 11220 9824
rect 11156 9764 11160 9820
rect 11160 9764 11216 9820
rect 11216 9764 11220 9820
rect 11156 9760 11220 9764
rect 11236 9820 11300 9824
rect 11236 9764 11240 9820
rect 11240 9764 11296 9820
rect 11296 9764 11300 9820
rect 11236 9760 11300 9764
rect 16916 9820 16980 9824
rect 16916 9764 16920 9820
rect 16920 9764 16976 9820
rect 16976 9764 16980 9820
rect 16916 9760 16980 9764
rect 16996 9820 17060 9824
rect 16996 9764 17000 9820
rect 17000 9764 17056 9820
rect 17056 9764 17060 9820
rect 16996 9760 17060 9764
rect 17076 9820 17140 9824
rect 17076 9764 17080 9820
rect 17080 9764 17136 9820
rect 17136 9764 17140 9820
rect 17076 9760 17140 9764
rect 17156 9820 17220 9824
rect 17156 9764 17160 9820
rect 17160 9764 17216 9820
rect 17216 9764 17220 9820
rect 17156 9760 17220 9764
rect 17236 9820 17300 9824
rect 17236 9764 17240 9820
rect 17240 9764 17296 9820
rect 17296 9764 17300 9820
rect 17236 9760 17300 9764
rect 22916 9820 22980 9824
rect 22916 9764 22920 9820
rect 22920 9764 22976 9820
rect 22976 9764 22980 9820
rect 22916 9760 22980 9764
rect 22996 9820 23060 9824
rect 22996 9764 23000 9820
rect 23000 9764 23056 9820
rect 23056 9764 23060 9820
rect 22996 9760 23060 9764
rect 23076 9820 23140 9824
rect 23076 9764 23080 9820
rect 23080 9764 23136 9820
rect 23136 9764 23140 9820
rect 23076 9760 23140 9764
rect 23156 9820 23220 9824
rect 23156 9764 23160 9820
rect 23160 9764 23216 9820
rect 23216 9764 23220 9820
rect 23156 9760 23220 9764
rect 23236 9820 23300 9824
rect 23236 9764 23240 9820
rect 23240 9764 23296 9820
rect 23296 9764 23300 9820
rect 23236 9760 23300 9764
rect 28916 9820 28980 9824
rect 28916 9764 28920 9820
rect 28920 9764 28976 9820
rect 28976 9764 28980 9820
rect 28916 9760 28980 9764
rect 28996 9820 29060 9824
rect 28996 9764 29000 9820
rect 29000 9764 29056 9820
rect 29056 9764 29060 9820
rect 28996 9760 29060 9764
rect 29076 9820 29140 9824
rect 29076 9764 29080 9820
rect 29080 9764 29136 9820
rect 29136 9764 29140 9820
rect 29076 9760 29140 9764
rect 29156 9820 29220 9824
rect 29156 9764 29160 9820
rect 29160 9764 29216 9820
rect 29216 9764 29220 9820
rect 29156 9760 29220 9764
rect 29236 9820 29300 9824
rect 29236 9764 29240 9820
rect 29240 9764 29296 9820
rect 29296 9764 29300 9820
rect 29236 9760 29300 9764
rect 4176 9276 4240 9280
rect 4176 9220 4180 9276
rect 4180 9220 4236 9276
rect 4236 9220 4240 9276
rect 4176 9216 4240 9220
rect 4256 9276 4320 9280
rect 4256 9220 4260 9276
rect 4260 9220 4316 9276
rect 4316 9220 4320 9276
rect 4256 9216 4320 9220
rect 4336 9276 4400 9280
rect 4336 9220 4340 9276
rect 4340 9220 4396 9276
rect 4396 9220 4400 9276
rect 4336 9216 4400 9220
rect 4416 9276 4480 9280
rect 4416 9220 4420 9276
rect 4420 9220 4476 9276
rect 4476 9220 4480 9276
rect 4416 9216 4480 9220
rect 4496 9276 4560 9280
rect 4496 9220 4500 9276
rect 4500 9220 4556 9276
rect 4556 9220 4560 9276
rect 4496 9216 4560 9220
rect 10176 9276 10240 9280
rect 10176 9220 10180 9276
rect 10180 9220 10236 9276
rect 10236 9220 10240 9276
rect 10176 9216 10240 9220
rect 10256 9276 10320 9280
rect 10256 9220 10260 9276
rect 10260 9220 10316 9276
rect 10316 9220 10320 9276
rect 10256 9216 10320 9220
rect 10336 9276 10400 9280
rect 10336 9220 10340 9276
rect 10340 9220 10396 9276
rect 10396 9220 10400 9276
rect 10336 9216 10400 9220
rect 10416 9276 10480 9280
rect 10416 9220 10420 9276
rect 10420 9220 10476 9276
rect 10476 9220 10480 9276
rect 10416 9216 10480 9220
rect 10496 9276 10560 9280
rect 10496 9220 10500 9276
rect 10500 9220 10556 9276
rect 10556 9220 10560 9276
rect 10496 9216 10560 9220
rect 16176 9276 16240 9280
rect 16176 9220 16180 9276
rect 16180 9220 16236 9276
rect 16236 9220 16240 9276
rect 16176 9216 16240 9220
rect 16256 9276 16320 9280
rect 16256 9220 16260 9276
rect 16260 9220 16316 9276
rect 16316 9220 16320 9276
rect 16256 9216 16320 9220
rect 16336 9276 16400 9280
rect 16336 9220 16340 9276
rect 16340 9220 16396 9276
rect 16396 9220 16400 9276
rect 16336 9216 16400 9220
rect 16416 9276 16480 9280
rect 16416 9220 16420 9276
rect 16420 9220 16476 9276
rect 16476 9220 16480 9276
rect 16416 9216 16480 9220
rect 16496 9276 16560 9280
rect 16496 9220 16500 9276
rect 16500 9220 16556 9276
rect 16556 9220 16560 9276
rect 16496 9216 16560 9220
rect 22176 9276 22240 9280
rect 22176 9220 22180 9276
rect 22180 9220 22236 9276
rect 22236 9220 22240 9276
rect 22176 9216 22240 9220
rect 22256 9276 22320 9280
rect 22256 9220 22260 9276
rect 22260 9220 22316 9276
rect 22316 9220 22320 9276
rect 22256 9216 22320 9220
rect 22336 9276 22400 9280
rect 22336 9220 22340 9276
rect 22340 9220 22396 9276
rect 22396 9220 22400 9276
rect 22336 9216 22400 9220
rect 22416 9276 22480 9280
rect 22416 9220 22420 9276
rect 22420 9220 22476 9276
rect 22476 9220 22480 9276
rect 22416 9216 22480 9220
rect 22496 9276 22560 9280
rect 22496 9220 22500 9276
rect 22500 9220 22556 9276
rect 22556 9220 22560 9276
rect 22496 9216 22560 9220
rect 28176 9276 28240 9280
rect 28176 9220 28180 9276
rect 28180 9220 28236 9276
rect 28236 9220 28240 9276
rect 28176 9216 28240 9220
rect 28256 9276 28320 9280
rect 28256 9220 28260 9276
rect 28260 9220 28316 9276
rect 28316 9220 28320 9276
rect 28256 9216 28320 9220
rect 28336 9276 28400 9280
rect 28336 9220 28340 9276
rect 28340 9220 28396 9276
rect 28396 9220 28400 9276
rect 28336 9216 28400 9220
rect 28416 9276 28480 9280
rect 28416 9220 28420 9276
rect 28420 9220 28476 9276
rect 28476 9220 28480 9276
rect 28416 9216 28480 9220
rect 28496 9276 28560 9280
rect 28496 9220 28500 9276
rect 28500 9220 28556 9276
rect 28556 9220 28560 9276
rect 28496 9216 28560 9220
rect 10732 8936 10796 8940
rect 10732 8880 10782 8936
rect 10782 8880 10796 8936
rect 10732 8876 10796 8880
rect 4916 8732 4980 8736
rect 4916 8676 4920 8732
rect 4920 8676 4976 8732
rect 4976 8676 4980 8732
rect 4916 8672 4980 8676
rect 4996 8732 5060 8736
rect 4996 8676 5000 8732
rect 5000 8676 5056 8732
rect 5056 8676 5060 8732
rect 4996 8672 5060 8676
rect 5076 8732 5140 8736
rect 5076 8676 5080 8732
rect 5080 8676 5136 8732
rect 5136 8676 5140 8732
rect 5076 8672 5140 8676
rect 5156 8732 5220 8736
rect 5156 8676 5160 8732
rect 5160 8676 5216 8732
rect 5216 8676 5220 8732
rect 5156 8672 5220 8676
rect 5236 8732 5300 8736
rect 5236 8676 5240 8732
rect 5240 8676 5296 8732
rect 5296 8676 5300 8732
rect 5236 8672 5300 8676
rect 10916 8732 10980 8736
rect 10916 8676 10920 8732
rect 10920 8676 10976 8732
rect 10976 8676 10980 8732
rect 10916 8672 10980 8676
rect 10996 8732 11060 8736
rect 10996 8676 11000 8732
rect 11000 8676 11056 8732
rect 11056 8676 11060 8732
rect 10996 8672 11060 8676
rect 11076 8732 11140 8736
rect 11076 8676 11080 8732
rect 11080 8676 11136 8732
rect 11136 8676 11140 8732
rect 11076 8672 11140 8676
rect 11156 8732 11220 8736
rect 11156 8676 11160 8732
rect 11160 8676 11216 8732
rect 11216 8676 11220 8732
rect 11156 8672 11220 8676
rect 11236 8732 11300 8736
rect 11236 8676 11240 8732
rect 11240 8676 11296 8732
rect 11296 8676 11300 8732
rect 11236 8672 11300 8676
rect 16916 8732 16980 8736
rect 16916 8676 16920 8732
rect 16920 8676 16976 8732
rect 16976 8676 16980 8732
rect 16916 8672 16980 8676
rect 16996 8732 17060 8736
rect 16996 8676 17000 8732
rect 17000 8676 17056 8732
rect 17056 8676 17060 8732
rect 16996 8672 17060 8676
rect 17076 8732 17140 8736
rect 17076 8676 17080 8732
rect 17080 8676 17136 8732
rect 17136 8676 17140 8732
rect 17076 8672 17140 8676
rect 17156 8732 17220 8736
rect 17156 8676 17160 8732
rect 17160 8676 17216 8732
rect 17216 8676 17220 8732
rect 17156 8672 17220 8676
rect 17236 8732 17300 8736
rect 17236 8676 17240 8732
rect 17240 8676 17296 8732
rect 17296 8676 17300 8732
rect 17236 8672 17300 8676
rect 22916 8732 22980 8736
rect 22916 8676 22920 8732
rect 22920 8676 22976 8732
rect 22976 8676 22980 8732
rect 22916 8672 22980 8676
rect 22996 8732 23060 8736
rect 22996 8676 23000 8732
rect 23000 8676 23056 8732
rect 23056 8676 23060 8732
rect 22996 8672 23060 8676
rect 23076 8732 23140 8736
rect 23076 8676 23080 8732
rect 23080 8676 23136 8732
rect 23136 8676 23140 8732
rect 23076 8672 23140 8676
rect 23156 8732 23220 8736
rect 23156 8676 23160 8732
rect 23160 8676 23216 8732
rect 23216 8676 23220 8732
rect 23156 8672 23220 8676
rect 23236 8732 23300 8736
rect 23236 8676 23240 8732
rect 23240 8676 23296 8732
rect 23296 8676 23300 8732
rect 23236 8672 23300 8676
rect 28916 8732 28980 8736
rect 28916 8676 28920 8732
rect 28920 8676 28976 8732
rect 28976 8676 28980 8732
rect 28916 8672 28980 8676
rect 28996 8732 29060 8736
rect 28996 8676 29000 8732
rect 29000 8676 29056 8732
rect 29056 8676 29060 8732
rect 28996 8672 29060 8676
rect 29076 8732 29140 8736
rect 29076 8676 29080 8732
rect 29080 8676 29136 8732
rect 29136 8676 29140 8732
rect 29076 8672 29140 8676
rect 29156 8732 29220 8736
rect 29156 8676 29160 8732
rect 29160 8676 29216 8732
rect 29216 8676 29220 8732
rect 29156 8672 29220 8676
rect 29236 8732 29300 8736
rect 29236 8676 29240 8732
rect 29240 8676 29296 8732
rect 29296 8676 29300 8732
rect 29236 8672 29300 8676
rect 9996 8528 10060 8532
rect 9996 8472 10046 8528
rect 10046 8472 10060 8528
rect 9996 8468 10060 8472
rect 4176 8188 4240 8192
rect 4176 8132 4180 8188
rect 4180 8132 4236 8188
rect 4236 8132 4240 8188
rect 4176 8128 4240 8132
rect 4256 8188 4320 8192
rect 4256 8132 4260 8188
rect 4260 8132 4316 8188
rect 4316 8132 4320 8188
rect 4256 8128 4320 8132
rect 4336 8188 4400 8192
rect 4336 8132 4340 8188
rect 4340 8132 4396 8188
rect 4396 8132 4400 8188
rect 4336 8128 4400 8132
rect 4416 8188 4480 8192
rect 4416 8132 4420 8188
rect 4420 8132 4476 8188
rect 4476 8132 4480 8188
rect 4416 8128 4480 8132
rect 4496 8188 4560 8192
rect 4496 8132 4500 8188
rect 4500 8132 4556 8188
rect 4556 8132 4560 8188
rect 4496 8128 4560 8132
rect 10176 8188 10240 8192
rect 10176 8132 10180 8188
rect 10180 8132 10236 8188
rect 10236 8132 10240 8188
rect 10176 8128 10240 8132
rect 10256 8188 10320 8192
rect 10256 8132 10260 8188
rect 10260 8132 10316 8188
rect 10316 8132 10320 8188
rect 10256 8128 10320 8132
rect 10336 8188 10400 8192
rect 10336 8132 10340 8188
rect 10340 8132 10396 8188
rect 10396 8132 10400 8188
rect 10336 8128 10400 8132
rect 10416 8188 10480 8192
rect 10416 8132 10420 8188
rect 10420 8132 10476 8188
rect 10476 8132 10480 8188
rect 10416 8128 10480 8132
rect 10496 8188 10560 8192
rect 10496 8132 10500 8188
rect 10500 8132 10556 8188
rect 10556 8132 10560 8188
rect 10496 8128 10560 8132
rect 16176 8188 16240 8192
rect 16176 8132 16180 8188
rect 16180 8132 16236 8188
rect 16236 8132 16240 8188
rect 16176 8128 16240 8132
rect 16256 8188 16320 8192
rect 16256 8132 16260 8188
rect 16260 8132 16316 8188
rect 16316 8132 16320 8188
rect 16256 8128 16320 8132
rect 16336 8188 16400 8192
rect 16336 8132 16340 8188
rect 16340 8132 16396 8188
rect 16396 8132 16400 8188
rect 16336 8128 16400 8132
rect 16416 8188 16480 8192
rect 16416 8132 16420 8188
rect 16420 8132 16476 8188
rect 16476 8132 16480 8188
rect 16416 8128 16480 8132
rect 16496 8188 16560 8192
rect 16496 8132 16500 8188
rect 16500 8132 16556 8188
rect 16556 8132 16560 8188
rect 16496 8128 16560 8132
rect 22176 8188 22240 8192
rect 22176 8132 22180 8188
rect 22180 8132 22236 8188
rect 22236 8132 22240 8188
rect 22176 8128 22240 8132
rect 22256 8188 22320 8192
rect 22256 8132 22260 8188
rect 22260 8132 22316 8188
rect 22316 8132 22320 8188
rect 22256 8128 22320 8132
rect 22336 8188 22400 8192
rect 22336 8132 22340 8188
rect 22340 8132 22396 8188
rect 22396 8132 22400 8188
rect 22336 8128 22400 8132
rect 22416 8188 22480 8192
rect 22416 8132 22420 8188
rect 22420 8132 22476 8188
rect 22476 8132 22480 8188
rect 22416 8128 22480 8132
rect 22496 8188 22560 8192
rect 22496 8132 22500 8188
rect 22500 8132 22556 8188
rect 22556 8132 22560 8188
rect 22496 8128 22560 8132
rect 28176 8188 28240 8192
rect 28176 8132 28180 8188
rect 28180 8132 28236 8188
rect 28236 8132 28240 8188
rect 28176 8128 28240 8132
rect 28256 8188 28320 8192
rect 28256 8132 28260 8188
rect 28260 8132 28316 8188
rect 28316 8132 28320 8188
rect 28256 8128 28320 8132
rect 28336 8188 28400 8192
rect 28336 8132 28340 8188
rect 28340 8132 28396 8188
rect 28396 8132 28400 8188
rect 28336 8128 28400 8132
rect 28416 8188 28480 8192
rect 28416 8132 28420 8188
rect 28420 8132 28476 8188
rect 28476 8132 28480 8188
rect 28416 8128 28480 8132
rect 28496 8188 28560 8192
rect 28496 8132 28500 8188
rect 28500 8132 28556 8188
rect 28556 8132 28560 8188
rect 28496 8128 28560 8132
rect 4916 7644 4980 7648
rect 4916 7588 4920 7644
rect 4920 7588 4976 7644
rect 4976 7588 4980 7644
rect 4916 7584 4980 7588
rect 4996 7644 5060 7648
rect 4996 7588 5000 7644
rect 5000 7588 5056 7644
rect 5056 7588 5060 7644
rect 4996 7584 5060 7588
rect 5076 7644 5140 7648
rect 5076 7588 5080 7644
rect 5080 7588 5136 7644
rect 5136 7588 5140 7644
rect 5076 7584 5140 7588
rect 5156 7644 5220 7648
rect 5156 7588 5160 7644
rect 5160 7588 5216 7644
rect 5216 7588 5220 7644
rect 5156 7584 5220 7588
rect 5236 7644 5300 7648
rect 5236 7588 5240 7644
rect 5240 7588 5296 7644
rect 5296 7588 5300 7644
rect 5236 7584 5300 7588
rect 10916 7644 10980 7648
rect 10916 7588 10920 7644
rect 10920 7588 10976 7644
rect 10976 7588 10980 7644
rect 10916 7584 10980 7588
rect 10996 7644 11060 7648
rect 10996 7588 11000 7644
rect 11000 7588 11056 7644
rect 11056 7588 11060 7644
rect 10996 7584 11060 7588
rect 11076 7644 11140 7648
rect 11076 7588 11080 7644
rect 11080 7588 11136 7644
rect 11136 7588 11140 7644
rect 11076 7584 11140 7588
rect 11156 7644 11220 7648
rect 11156 7588 11160 7644
rect 11160 7588 11216 7644
rect 11216 7588 11220 7644
rect 11156 7584 11220 7588
rect 11236 7644 11300 7648
rect 11236 7588 11240 7644
rect 11240 7588 11296 7644
rect 11296 7588 11300 7644
rect 11236 7584 11300 7588
rect 16916 7644 16980 7648
rect 16916 7588 16920 7644
rect 16920 7588 16976 7644
rect 16976 7588 16980 7644
rect 16916 7584 16980 7588
rect 16996 7644 17060 7648
rect 16996 7588 17000 7644
rect 17000 7588 17056 7644
rect 17056 7588 17060 7644
rect 16996 7584 17060 7588
rect 17076 7644 17140 7648
rect 17076 7588 17080 7644
rect 17080 7588 17136 7644
rect 17136 7588 17140 7644
rect 17076 7584 17140 7588
rect 17156 7644 17220 7648
rect 17156 7588 17160 7644
rect 17160 7588 17216 7644
rect 17216 7588 17220 7644
rect 17156 7584 17220 7588
rect 17236 7644 17300 7648
rect 17236 7588 17240 7644
rect 17240 7588 17296 7644
rect 17296 7588 17300 7644
rect 17236 7584 17300 7588
rect 22916 7644 22980 7648
rect 22916 7588 22920 7644
rect 22920 7588 22976 7644
rect 22976 7588 22980 7644
rect 22916 7584 22980 7588
rect 22996 7644 23060 7648
rect 22996 7588 23000 7644
rect 23000 7588 23056 7644
rect 23056 7588 23060 7644
rect 22996 7584 23060 7588
rect 23076 7644 23140 7648
rect 23076 7588 23080 7644
rect 23080 7588 23136 7644
rect 23136 7588 23140 7644
rect 23076 7584 23140 7588
rect 23156 7644 23220 7648
rect 23156 7588 23160 7644
rect 23160 7588 23216 7644
rect 23216 7588 23220 7644
rect 23156 7584 23220 7588
rect 23236 7644 23300 7648
rect 23236 7588 23240 7644
rect 23240 7588 23296 7644
rect 23296 7588 23300 7644
rect 23236 7584 23300 7588
rect 28916 7644 28980 7648
rect 28916 7588 28920 7644
rect 28920 7588 28976 7644
rect 28976 7588 28980 7644
rect 28916 7584 28980 7588
rect 28996 7644 29060 7648
rect 28996 7588 29000 7644
rect 29000 7588 29056 7644
rect 29056 7588 29060 7644
rect 28996 7584 29060 7588
rect 29076 7644 29140 7648
rect 29076 7588 29080 7644
rect 29080 7588 29136 7644
rect 29136 7588 29140 7644
rect 29076 7584 29140 7588
rect 29156 7644 29220 7648
rect 29156 7588 29160 7644
rect 29160 7588 29216 7644
rect 29216 7588 29220 7644
rect 29156 7584 29220 7588
rect 29236 7644 29300 7648
rect 29236 7588 29240 7644
rect 29240 7588 29296 7644
rect 29296 7588 29300 7644
rect 29236 7584 29300 7588
rect 4176 7100 4240 7104
rect 4176 7044 4180 7100
rect 4180 7044 4236 7100
rect 4236 7044 4240 7100
rect 4176 7040 4240 7044
rect 4256 7100 4320 7104
rect 4256 7044 4260 7100
rect 4260 7044 4316 7100
rect 4316 7044 4320 7100
rect 4256 7040 4320 7044
rect 4336 7100 4400 7104
rect 4336 7044 4340 7100
rect 4340 7044 4396 7100
rect 4396 7044 4400 7100
rect 4336 7040 4400 7044
rect 4416 7100 4480 7104
rect 4416 7044 4420 7100
rect 4420 7044 4476 7100
rect 4476 7044 4480 7100
rect 4416 7040 4480 7044
rect 4496 7100 4560 7104
rect 4496 7044 4500 7100
rect 4500 7044 4556 7100
rect 4556 7044 4560 7100
rect 4496 7040 4560 7044
rect 10176 7100 10240 7104
rect 10176 7044 10180 7100
rect 10180 7044 10236 7100
rect 10236 7044 10240 7100
rect 10176 7040 10240 7044
rect 10256 7100 10320 7104
rect 10256 7044 10260 7100
rect 10260 7044 10316 7100
rect 10316 7044 10320 7100
rect 10256 7040 10320 7044
rect 10336 7100 10400 7104
rect 10336 7044 10340 7100
rect 10340 7044 10396 7100
rect 10396 7044 10400 7100
rect 10336 7040 10400 7044
rect 10416 7100 10480 7104
rect 10416 7044 10420 7100
rect 10420 7044 10476 7100
rect 10476 7044 10480 7100
rect 10416 7040 10480 7044
rect 10496 7100 10560 7104
rect 10496 7044 10500 7100
rect 10500 7044 10556 7100
rect 10556 7044 10560 7100
rect 10496 7040 10560 7044
rect 16176 7100 16240 7104
rect 16176 7044 16180 7100
rect 16180 7044 16236 7100
rect 16236 7044 16240 7100
rect 16176 7040 16240 7044
rect 16256 7100 16320 7104
rect 16256 7044 16260 7100
rect 16260 7044 16316 7100
rect 16316 7044 16320 7100
rect 16256 7040 16320 7044
rect 16336 7100 16400 7104
rect 16336 7044 16340 7100
rect 16340 7044 16396 7100
rect 16396 7044 16400 7100
rect 16336 7040 16400 7044
rect 16416 7100 16480 7104
rect 16416 7044 16420 7100
rect 16420 7044 16476 7100
rect 16476 7044 16480 7100
rect 16416 7040 16480 7044
rect 16496 7100 16560 7104
rect 16496 7044 16500 7100
rect 16500 7044 16556 7100
rect 16556 7044 16560 7100
rect 16496 7040 16560 7044
rect 22176 7100 22240 7104
rect 22176 7044 22180 7100
rect 22180 7044 22236 7100
rect 22236 7044 22240 7100
rect 22176 7040 22240 7044
rect 22256 7100 22320 7104
rect 22256 7044 22260 7100
rect 22260 7044 22316 7100
rect 22316 7044 22320 7100
rect 22256 7040 22320 7044
rect 22336 7100 22400 7104
rect 22336 7044 22340 7100
rect 22340 7044 22396 7100
rect 22396 7044 22400 7100
rect 22336 7040 22400 7044
rect 22416 7100 22480 7104
rect 22416 7044 22420 7100
rect 22420 7044 22476 7100
rect 22476 7044 22480 7100
rect 22416 7040 22480 7044
rect 22496 7100 22560 7104
rect 22496 7044 22500 7100
rect 22500 7044 22556 7100
rect 22556 7044 22560 7100
rect 22496 7040 22560 7044
rect 28176 7100 28240 7104
rect 28176 7044 28180 7100
rect 28180 7044 28236 7100
rect 28236 7044 28240 7100
rect 28176 7040 28240 7044
rect 28256 7100 28320 7104
rect 28256 7044 28260 7100
rect 28260 7044 28316 7100
rect 28316 7044 28320 7100
rect 28256 7040 28320 7044
rect 28336 7100 28400 7104
rect 28336 7044 28340 7100
rect 28340 7044 28396 7100
rect 28396 7044 28400 7100
rect 28336 7040 28400 7044
rect 28416 7100 28480 7104
rect 28416 7044 28420 7100
rect 28420 7044 28476 7100
rect 28476 7044 28480 7100
rect 28416 7040 28480 7044
rect 28496 7100 28560 7104
rect 28496 7044 28500 7100
rect 28500 7044 28556 7100
rect 28556 7044 28560 7100
rect 28496 7040 28560 7044
rect 10732 6700 10796 6764
rect 4916 6556 4980 6560
rect 4916 6500 4920 6556
rect 4920 6500 4976 6556
rect 4976 6500 4980 6556
rect 4916 6496 4980 6500
rect 4996 6556 5060 6560
rect 4996 6500 5000 6556
rect 5000 6500 5056 6556
rect 5056 6500 5060 6556
rect 4996 6496 5060 6500
rect 5076 6556 5140 6560
rect 5076 6500 5080 6556
rect 5080 6500 5136 6556
rect 5136 6500 5140 6556
rect 5076 6496 5140 6500
rect 5156 6556 5220 6560
rect 5156 6500 5160 6556
rect 5160 6500 5216 6556
rect 5216 6500 5220 6556
rect 5156 6496 5220 6500
rect 5236 6556 5300 6560
rect 5236 6500 5240 6556
rect 5240 6500 5296 6556
rect 5296 6500 5300 6556
rect 5236 6496 5300 6500
rect 10916 6556 10980 6560
rect 10916 6500 10920 6556
rect 10920 6500 10976 6556
rect 10976 6500 10980 6556
rect 10916 6496 10980 6500
rect 10996 6556 11060 6560
rect 10996 6500 11000 6556
rect 11000 6500 11056 6556
rect 11056 6500 11060 6556
rect 10996 6496 11060 6500
rect 11076 6556 11140 6560
rect 11076 6500 11080 6556
rect 11080 6500 11136 6556
rect 11136 6500 11140 6556
rect 11076 6496 11140 6500
rect 11156 6556 11220 6560
rect 11156 6500 11160 6556
rect 11160 6500 11216 6556
rect 11216 6500 11220 6556
rect 11156 6496 11220 6500
rect 11236 6556 11300 6560
rect 11236 6500 11240 6556
rect 11240 6500 11296 6556
rect 11296 6500 11300 6556
rect 11236 6496 11300 6500
rect 16916 6556 16980 6560
rect 16916 6500 16920 6556
rect 16920 6500 16976 6556
rect 16976 6500 16980 6556
rect 16916 6496 16980 6500
rect 16996 6556 17060 6560
rect 16996 6500 17000 6556
rect 17000 6500 17056 6556
rect 17056 6500 17060 6556
rect 16996 6496 17060 6500
rect 17076 6556 17140 6560
rect 17076 6500 17080 6556
rect 17080 6500 17136 6556
rect 17136 6500 17140 6556
rect 17076 6496 17140 6500
rect 17156 6556 17220 6560
rect 17156 6500 17160 6556
rect 17160 6500 17216 6556
rect 17216 6500 17220 6556
rect 17156 6496 17220 6500
rect 17236 6556 17300 6560
rect 17236 6500 17240 6556
rect 17240 6500 17296 6556
rect 17296 6500 17300 6556
rect 17236 6496 17300 6500
rect 22916 6556 22980 6560
rect 22916 6500 22920 6556
rect 22920 6500 22976 6556
rect 22976 6500 22980 6556
rect 22916 6496 22980 6500
rect 22996 6556 23060 6560
rect 22996 6500 23000 6556
rect 23000 6500 23056 6556
rect 23056 6500 23060 6556
rect 22996 6496 23060 6500
rect 23076 6556 23140 6560
rect 23076 6500 23080 6556
rect 23080 6500 23136 6556
rect 23136 6500 23140 6556
rect 23076 6496 23140 6500
rect 23156 6556 23220 6560
rect 23156 6500 23160 6556
rect 23160 6500 23216 6556
rect 23216 6500 23220 6556
rect 23156 6496 23220 6500
rect 23236 6556 23300 6560
rect 23236 6500 23240 6556
rect 23240 6500 23296 6556
rect 23296 6500 23300 6556
rect 23236 6496 23300 6500
rect 28916 6556 28980 6560
rect 28916 6500 28920 6556
rect 28920 6500 28976 6556
rect 28976 6500 28980 6556
rect 28916 6496 28980 6500
rect 28996 6556 29060 6560
rect 28996 6500 29000 6556
rect 29000 6500 29056 6556
rect 29056 6500 29060 6556
rect 28996 6496 29060 6500
rect 29076 6556 29140 6560
rect 29076 6500 29080 6556
rect 29080 6500 29136 6556
rect 29136 6500 29140 6556
rect 29076 6496 29140 6500
rect 29156 6556 29220 6560
rect 29156 6500 29160 6556
rect 29160 6500 29216 6556
rect 29216 6500 29220 6556
rect 29156 6496 29220 6500
rect 29236 6556 29300 6560
rect 29236 6500 29240 6556
rect 29240 6500 29296 6556
rect 29296 6500 29300 6556
rect 29236 6496 29300 6500
rect 4176 6012 4240 6016
rect 4176 5956 4180 6012
rect 4180 5956 4236 6012
rect 4236 5956 4240 6012
rect 4176 5952 4240 5956
rect 4256 6012 4320 6016
rect 4256 5956 4260 6012
rect 4260 5956 4316 6012
rect 4316 5956 4320 6012
rect 4256 5952 4320 5956
rect 4336 6012 4400 6016
rect 4336 5956 4340 6012
rect 4340 5956 4396 6012
rect 4396 5956 4400 6012
rect 4336 5952 4400 5956
rect 4416 6012 4480 6016
rect 4416 5956 4420 6012
rect 4420 5956 4476 6012
rect 4476 5956 4480 6012
rect 4416 5952 4480 5956
rect 4496 6012 4560 6016
rect 4496 5956 4500 6012
rect 4500 5956 4556 6012
rect 4556 5956 4560 6012
rect 4496 5952 4560 5956
rect 10176 6012 10240 6016
rect 10176 5956 10180 6012
rect 10180 5956 10236 6012
rect 10236 5956 10240 6012
rect 10176 5952 10240 5956
rect 10256 6012 10320 6016
rect 10256 5956 10260 6012
rect 10260 5956 10316 6012
rect 10316 5956 10320 6012
rect 10256 5952 10320 5956
rect 10336 6012 10400 6016
rect 10336 5956 10340 6012
rect 10340 5956 10396 6012
rect 10396 5956 10400 6012
rect 10336 5952 10400 5956
rect 10416 6012 10480 6016
rect 10416 5956 10420 6012
rect 10420 5956 10476 6012
rect 10476 5956 10480 6012
rect 10416 5952 10480 5956
rect 10496 6012 10560 6016
rect 10496 5956 10500 6012
rect 10500 5956 10556 6012
rect 10556 5956 10560 6012
rect 10496 5952 10560 5956
rect 16176 6012 16240 6016
rect 16176 5956 16180 6012
rect 16180 5956 16236 6012
rect 16236 5956 16240 6012
rect 16176 5952 16240 5956
rect 16256 6012 16320 6016
rect 16256 5956 16260 6012
rect 16260 5956 16316 6012
rect 16316 5956 16320 6012
rect 16256 5952 16320 5956
rect 16336 6012 16400 6016
rect 16336 5956 16340 6012
rect 16340 5956 16396 6012
rect 16396 5956 16400 6012
rect 16336 5952 16400 5956
rect 16416 6012 16480 6016
rect 16416 5956 16420 6012
rect 16420 5956 16476 6012
rect 16476 5956 16480 6012
rect 16416 5952 16480 5956
rect 16496 6012 16560 6016
rect 16496 5956 16500 6012
rect 16500 5956 16556 6012
rect 16556 5956 16560 6012
rect 16496 5952 16560 5956
rect 22176 6012 22240 6016
rect 22176 5956 22180 6012
rect 22180 5956 22236 6012
rect 22236 5956 22240 6012
rect 22176 5952 22240 5956
rect 22256 6012 22320 6016
rect 22256 5956 22260 6012
rect 22260 5956 22316 6012
rect 22316 5956 22320 6012
rect 22256 5952 22320 5956
rect 22336 6012 22400 6016
rect 22336 5956 22340 6012
rect 22340 5956 22396 6012
rect 22396 5956 22400 6012
rect 22336 5952 22400 5956
rect 22416 6012 22480 6016
rect 22416 5956 22420 6012
rect 22420 5956 22476 6012
rect 22476 5956 22480 6012
rect 22416 5952 22480 5956
rect 22496 6012 22560 6016
rect 22496 5956 22500 6012
rect 22500 5956 22556 6012
rect 22556 5956 22560 6012
rect 22496 5952 22560 5956
rect 28176 6012 28240 6016
rect 28176 5956 28180 6012
rect 28180 5956 28236 6012
rect 28236 5956 28240 6012
rect 28176 5952 28240 5956
rect 28256 6012 28320 6016
rect 28256 5956 28260 6012
rect 28260 5956 28316 6012
rect 28316 5956 28320 6012
rect 28256 5952 28320 5956
rect 28336 6012 28400 6016
rect 28336 5956 28340 6012
rect 28340 5956 28396 6012
rect 28396 5956 28400 6012
rect 28336 5952 28400 5956
rect 28416 6012 28480 6016
rect 28416 5956 28420 6012
rect 28420 5956 28476 6012
rect 28476 5956 28480 6012
rect 28416 5952 28480 5956
rect 28496 6012 28560 6016
rect 28496 5956 28500 6012
rect 28500 5956 28556 6012
rect 28556 5956 28560 6012
rect 28496 5952 28560 5956
rect 4916 5468 4980 5472
rect 4916 5412 4920 5468
rect 4920 5412 4976 5468
rect 4976 5412 4980 5468
rect 4916 5408 4980 5412
rect 4996 5468 5060 5472
rect 4996 5412 5000 5468
rect 5000 5412 5056 5468
rect 5056 5412 5060 5468
rect 4996 5408 5060 5412
rect 5076 5468 5140 5472
rect 5076 5412 5080 5468
rect 5080 5412 5136 5468
rect 5136 5412 5140 5468
rect 5076 5408 5140 5412
rect 5156 5468 5220 5472
rect 5156 5412 5160 5468
rect 5160 5412 5216 5468
rect 5216 5412 5220 5468
rect 5156 5408 5220 5412
rect 5236 5468 5300 5472
rect 5236 5412 5240 5468
rect 5240 5412 5296 5468
rect 5296 5412 5300 5468
rect 5236 5408 5300 5412
rect 10916 5468 10980 5472
rect 10916 5412 10920 5468
rect 10920 5412 10976 5468
rect 10976 5412 10980 5468
rect 10916 5408 10980 5412
rect 10996 5468 11060 5472
rect 10996 5412 11000 5468
rect 11000 5412 11056 5468
rect 11056 5412 11060 5468
rect 10996 5408 11060 5412
rect 11076 5468 11140 5472
rect 11076 5412 11080 5468
rect 11080 5412 11136 5468
rect 11136 5412 11140 5468
rect 11076 5408 11140 5412
rect 11156 5468 11220 5472
rect 11156 5412 11160 5468
rect 11160 5412 11216 5468
rect 11216 5412 11220 5468
rect 11156 5408 11220 5412
rect 11236 5468 11300 5472
rect 11236 5412 11240 5468
rect 11240 5412 11296 5468
rect 11296 5412 11300 5468
rect 11236 5408 11300 5412
rect 16916 5468 16980 5472
rect 16916 5412 16920 5468
rect 16920 5412 16976 5468
rect 16976 5412 16980 5468
rect 16916 5408 16980 5412
rect 16996 5468 17060 5472
rect 16996 5412 17000 5468
rect 17000 5412 17056 5468
rect 17056 5412 17060 5468
rect 16996 5408 17060 5412
rect 17076 5468 17140 5472
rect 17076 5412 17080 5468
rect 17080 5412 17136 5468
rect 17136 5412 17140 5468
rect 17076 5408 17140 5412
rect 17156 5468 17220 5472
rect 17156 5412 17160 5468
rect 17160 5412 17216 5468
rect 17216 5412 17220 5468
rect 17156 5408 17220 5412
rect 17236 5468 17300 5472
rect 17236 5412 17240 5468
rect 17240 5412 17296 5468
rect 17296 5412 17300 5468
rect 17236 5408 17300 5412
rect 22916 5468 22980 5472
rect 22916 5412 22920 5468
rect 22920 5412 22976 5468
rect 22976 5412 22980 5468
rect 22916 5408 22980 5412
rect 22996 5468 23060 5472
rect 22996 5412 23000 5468
rect 23000 5412 23056 5468
rect 23056 5412 23060 5468
rect 22996 5408 23060 5412
rect 23076 5468 23140 5472
rect 23076 5412 23080 5468
rect 23080 5412 23136 5468
rect 23136 5412 23140 5468
rect 23076 5408 23140 5412
rect 23156 5468 23220 5472
rect 23156 5412 23160 5468
rect 23160 5412 23216 5468
rect 23216 5412 23220 5468
rect 23156 5408 23220 5412
rect 23236 5468 23300 5472
rect 23236 5412 23240 5468
rect 23240 5412 23296 5468
rect 23296 5412 23300 5468
rect 23236 5408 23300 5412
rect 28916 5468 28980 5472
rect 28916 5412 28920 5468
rect 28920 5412 28976 5468
rect 28976 5412 28980 5468
rect 28916 5408 28980 5412
rect 28996 5468 29060 5472
rect 28996 5412 29000 5468
rect 29000 5412 29056 5468
rect 29056 5412 29060 5468
rect 28996 5408 29060 5412
rect 29076 5468 29140 5472
rect 29076 5412 29080 5468
rect 29080 5412 29136 5468
rect 29136 5412 29140 5468
rect 29076 5408 29140 5412
rect 29156 5468 29220 5472
rect 29156 5412 29160 5468
rect 29160 5412 29216 5468
rect 29216 5412 29220 5468
rect 29156 5408 29220 5412
rect 29236 5468 29300 5472
rect 29236 5412 29240 5468
rect 29240 5412 29296 5468
rect 29296 5412 29300 5468
rect 29236 5408 29300 5412
rect 9996 4992 10060 4996
rect 9996 4936 10046 4992
rect 10046 4936 10060 4992
rect 9996 4932 10060 4936
rect 4176 4924 4240 4928
rect 4176 4868 4180 4924
rect 4180 4868 4236 4924
rect 4236 4868 4240 4924
rect 4176 4864 4240 4868
rect 4256 4924 4320 4928
rect 4256 4868 4260 4924
rect 4260 4868 4316 4924
rect 4316 4868 4320 4924
rect 4256 4864 4320 4868
rect 4336 4924 4400 4928
rect 4336 4868 4340 4924
rect 4340 4868 4396 4924
rect 4396 4868 4400 4924
rect 4336 4864 4400 4868
rect 4416 4924 4480 4928
rect 4416 4868 4420 4924
rect 4420 4868 4476 4924
rect 4476 4868 4480 4924
rect 4416 4864 4480 4868
rect 4496 4924 4560 4928
rect 4496 4868 4500 4924
rect 4500 4868 4556 4924
rect 4556 4868 4560 4924
rect 4496 4864 4560 4868
rect 10176 4924 10240 4928
rect 10176 4868 10180 4924
rect 10180 4868 10236 4924
rect 10236 4868 10240 4924
rect 10176 4864 10240 4868
rect 10256 4924 10320 4928
rect 10256 4868 10260 4924
rect 10260 4868 10316 4924
rect 10316 4868 10320 4924
rect 10256 4864 10320 4868
rect 10336 4924 10400 4928
rect 10336 4868 10340 4924
rect 10340 4868 10396 4924
rect 10396 4868 10400 4924
rect 10336 4864 10400 4868
rect 10416 4924 10480 4928
rect 10416 4868 10420 4924
rect 10420 4868 10476 4924
rect 10476 4868 10480 4924
rect 10416 4864 10480 4868
rect 10496 4924 10560 4928
rect 10496 4868 10500 4924
rect 10500 4868 10556 4924
rect 10556 4868 10560 4924
rect 10496 4864 10560 4868
rect 16176 4924 16240 4928
rect 16176 4868 16180 4924
rect 16180 4868 16236 4924
rect 16236 4868 16240 4924
rect 16176 4864 16240 4868
rect 16256 4924 16320 4928
rect 16256 4868 16260 4924
rect 16260 4868 16316 4924
rect 16316 4868 16320 4924
rect 16256 4864 16320 4868
rect 16336 4924 16400 4928
rect 16336 4868 16340 4924
rect 16340 4868 16396 4924
rect 16396 4868 16400 4924
rect 16336 4864 16400 4868
rect 16416 4924 16480 4928
rect 16416 4868 16420 4924
rect 16420 4868 16476 4924
rect 16476 4868 16480 4924
rect 16416 4864 16480 4868
rect 16496 4924 16560 4928
rect 16496 4868 16500 4924
rect 16500 4868 16556 4924
rect 16556 4868 16560 4924
rect 16496 4864 16560 4868
rect 22176 4924 22240 4928
rect 22176 4868 22180 4924
rect 22180 4868 22236 4924
rect 22236 4868 22240 4924
rect 22176 4864 22240 4868
rect 22256 4924 22320 4928
rect 22256 4868 22260 4924
rect 22260 4868 22316 4924
rect 22316 4868 22320 4924
rect 22256 4864 22320 4868
rect 22336 4924 22400 4928
rect 22336 4868 22340 4924
rect 22340 4868 22396 4924
rect 22396 4868 22400 4924
rect 22336 4864 22400 4868
rect 22416 4924 22480 4928
rect 22416 4868 22420 4924
rect 22420 4868 22476 4924
rect 22476 4868 22480 4924
rect 22416 4864 22480 4868
rect 22496 4924 22560 4928
rect 22496 4868 22500 4924
rect 22500 4868 22556 4924
rect 22556 4868 22560 4924
rect 22496 4864 22560 4868
rect 28176 4924 28240 4928
rect 28176 4868 28180 4924
rect 28180 4868 28236 4924
rect 28236 4868 28240 4924
rect 28176 4864 28240 4868
rect 28256 4924 28320 4928
rect 28256 4868 28260 4924
rect 28260 4868 28316 4924
rect 28316 4868 28320 4924
rect 28256 4864 28320 4868
rect 28336 4924 28400 4928
rect 28336 4868 28340 4924
rect 28340 4868 28396 4924
rect 28396 4868 28400 4924
rect 28336 4864 28400 4868
rect 28416 4924 28480 4928
rect 28416 4868 28420 4924
rect 28420 4868 28476 4924
rect 28476 4868 28480 4924
rect 28416 4864 28480 4868
rect 28496 4924 28560 4928
rect 28496 4868 28500 4924
rect 28500 4868 28556 4924
rect 28556 4868 28560 4924
rect 28496 4864 28560 4868
rect 4916 4380 4980 4384
rect 4916 4324 4920 4380
rect 4920 4324 4976 4380
rect 4976 4324 4980 4380
rect 4916 4320 4980 4324
rect 4996 4380 5060 4384
rect 4996 4324 5000 4380
rect 5000 4324 5056 4380
rect 5056 4324 5060 4380
rect 4996 4320 5060 4324
rect 5076 4380 5140 4384
rect 5076 4324 5080 4380
rect 5080 4324 5136 4380
rect 5136 4324 5140 4380
rect 5076 4320 5140 4324
rect 5156 4380 5220 4384
rect 5156 4324 5160 4380
rect 5160 4324 5216 4380
rect 5216 4324 5220 4380
rect 5156 4320 5220 4324
rect 5236 4380 5300 4384
rect 5236 4324 5240 4380
rect 5240 4324 5296 4380
rect 5296 4324 5300 4380
rect 5236 4320 5300 4324
rect 10916 4380 10980 4384
rect 10916 4324 10920 4380
rect 10920 4324 10976 4380
rect 10976 4324 10980 4380
rect 10916 4320 10980 4324
rect 10996 4380 11060 4384
rect 10996 4324 11000 4380
rect 11000 4324 11056 4380
rect 11056 4324 11060 4380
rect 10996 4320 11060 4324
rect 11076 4380 11140 4384
rect 11076 4324 11080 4380
rect 11080 4324 11136 4380
rect 11136 4324 11140 4380
rect 11076 4320 11140 4324
rect 11156 4380 11220 4384
rect 11156 4324 11160 4380
rect 11160 4324 11216 4380
rect 11216 4324 11220 4380
rect 11156 4320 11220 4324
rect 11236 4380 11300 4384
rect 11236 4324 11240 4380
rect 11240 4324 11296 4380
rect 11296 4324 11300 4380
rect 11236 4320 11300 4324
rect 16916 4380 16980 4384
rect 16916 4324 16920 4380
rect 16920 4324 16976 4380
rect 16976 4324 16980 4380
rect 16916 4320 16980 4324
rect 16996 4380 17060 4384
rect 16996 4324 17000 4380
rect 17000 4324 17056 4380
rect 17056 4324 17060 4380
rect 16996 4320 17060 4324
rect 17076 4380 17140 4384
rect 17076 4324 17080 4380
rect 17080 4324 17136 4380
rect 17136 4324 17140 4380
rect 17076 4320 17140 4324
rect 17156 4380 17220 4384
rect 17156 4324 17160 4380
rect 17160 4324 17216 4380
rect 17216 4324 17220 4380
rect 17156 4320 17220 4324
rect 17236 4380 17300 4384
rect 17236 4324 17240 4380
rect 17240 4324 17296 4380
rect 17296 4324 17300 4380
rect 17236 4320 17300 4324
rect 22916 4380 22980 4384
rect 22916 4324 22920 4380
rect 22920 4324 22976 4380
rect 22976 4324 22980 4380
rect 22916 4320 22980 4324
rect 22996 4380 23060 4384
rect 22996 4324 23000 4380
rect 23000 4324 23056 4380
rect 23056 4324 23060 4380
rect 22996 4320 23060 4324
rect 23076 4380 23140 4384
rect 23076 4324 23080 4380
rect 23080 4324 23136 4380
rect 23136 4324 23140 4380
rect 23076 4320 23140 4324
rect 23156 4380 23220 4384
rect 23156 4324 23160 4380
rect 23160 4324 23216 4380
rect 23216 4324 23220 4380
rect 23156 4320 23220 4324
rect 23236 4380 23300 4384
rect 23236 4324 23240 4380
rect 23240 4324 23296 4380
rect 23296 4324 23300 4380
rect 23236 4320 23300 4324
rect 28916 4380 28980 4384
rect 28916 4324 28920 4380
rect 28920 4324 28976 4380
rect 28976 4324 28980 4380
rect 28916 4320 28980 4324
rect 28996 4380 29060 4384
rect 28996 4324 29000 4380
rect 29000 4324 29056 4380
rect 29056 4324 29060 4380
rect 28996 4320 29060 4324
rect 29076 4380 29140 4384
rect 29076 4324 29080 4380
rect 29080 4324 29136 4380
rect 29136 4324 29140 4380
rect 29076 4320 29140 4324
rect 29156 4380 29220 4384
rect 29156 4324 29160 4380
rect 29160 4324 29216 4380
rect 29216 4324 29220 4380
rect 29156 4320 29220 4324
rect 29236 4380 29300 4384
rect 29236 4324 29240 4380
rect 29240 4324 29296 4380
rect 29296 4324 29300 4380
rect 29236 4320 29300 4324
rect 4176 3836 4240 3840
rect 4176 3780 4180 3836
rect 4180 3780 4236 3836
rect 4236 3780 4240 3836
rect 4176 3776 4240 3780
rect 4256 3836 4320 3840
rect 4256 3780 4260 3836
rect 4260 3780 4316 3836
rect 4316 3780 4320 3836
rect 4256 3776 4320 3780
rect 4336 3836 4400 3840
rect 4336 3780 4340 3836
rect 4340 3780 4396 3836
rect 4396 3780 4400 3836
rect 4336 3776 4400 3780
rect 4416 3836 4480 3840
rect 4416 3780 4420 3836
rect 4420 3780 4476 3836
rect 4476 3780 4480 3836
rect 4416 3776 4480 3780
rect 4496 3836 4560 3840
rect 4496 3780 4500 3836
rect 4500 3780 4556 3836
rect 4556 3780 4560 3836
rect 4496 3776 4560 3780
rect 10176 3836 10240 3840
rect 10176 3780 10180 3836
rect 10180 3780 10236 3836
rect 10236 3780 10240 3836
rect 10176 3776 10240 3780
rect 10256 3836 10320 3840
rect 10256 3780 10260 3836
rect 10260 3780 10316 3836
rect 10316 3780 10320 3836
rect 10256 3776 10320 3780
rect 10336 3836 10400 3840
rect 10336 3780 10340 3836
rect 10340 3780 10396 3836
rect 10396 3780 10400 3836
rect 10336 3776 10400 3780
rect 10416 3836 10480 3840
rect 10416 3780 10420 3836
rect 10420 3780 10476 3836
rect 10476 3780 10480 3836
rect 10416 3776 10480 3780
rect 10496 3836 10560 3840
rect 10496 3780 10500 3836
rect 10500 3780 10556 3836
rect 10556 3780 10560 3836
rect 10496 3776 10560 3780
rect 16176 3836 16240 3840
rect 16176 3780 16180 3836
rect 16180 3780 16236 3836
rect 16236 3780 16240 3836
rect 16176 3776 16240 3780
rect 16256 3836 16320 3840
rect 16256 3780 16260 3836
rect 16260 3780 16316 3836
rect 16316 3780 16320 3836
rect 16256 3776 16320 3780
rect 16336 3836 16400 3840
rect 16336 3780 16340 3836
rect 16340 3780 16396 3836
rect 16396 3780 16400 3836
rect 16336 3776 16400 3780
rect 16416 3836 16480 3840
rect 16416 3780 16420 3836
rect 16420 3780 16476 3836
rect 16476 3780 16480 3836
rect 16416 3776 16480 3780
rect 16496 3836 16560 3840
rect 16496 3780 16500 3836
rect 16500 3780 16556 3836
rect 16556 3780 16560 3836
rect 16496 3776 16560 3780
rect 22176 3836 22240 3840
rect 22176 3780 22180 3836
rect 22180 3780 22236 3836
rect 22236 3780 22240 3836
rect 22176 3776 22240 3780
rect 22256 3836 22320 3840
rect 22256 3780 22260 3836
rect 22260 3780 22316 3836
rect 22316 3780 22320 3836
rect 22256 3776 22320 3780
rect 22336 3836 22400 3840
rect 22336 3780 22340 3836
rect 22340 3780 22396 3836
rect 22396 3780 22400 3836
rect 22336 3776 22400 3780
rect 22416 3836 22480 3840
rect 22416 3780 22420 3836
rect 22420 3780 22476 3836
rect 22476 3780 22480 3836
rect 22416 3776 22480 3780
rect 22496 3836 22560 3840
rect 22496 3780 22500 3836
rect 22500 3780 22556 3836
rect 22556 3780 22560 3836
rect 22496 3776 22560 3780
rect 28176 3836 28240 3840
rect 28176 3780 28180 3836
rect 28180 3780 28236 3836
rect 28236 3780 28240 3836
rect 28176 3776 28240 3780
rect 28256 3836 28320 3840
rect 28256 3780 28260 3836
rect 28260 3780 28316 3836
rect 28316 3780 28320 3836
rect 28256 3776 28320 3780
rect 28336 3836 28400 3840
rect 28336 3780 28340 3836
rect 28340 3780 28396 3836
rect 28396 3780 28400 3836
rect 28336 3776 28400 3780
rect 28416 3836 28480 3840
rect 28416 3780 28420 3836
rect 28420 3780 28476 3836
rect 28476 3780 28480 3836
rect 28416 3776 28480 3780
rect 28496 3836 28560 3840
rect 28496 3780 28500 3836
rect 28500 3780 28556 3836
rect 28556 3780 28560 3836
rect 28496 3776 28560 3780
rect 4916 3292 4980 3296
rect 4916 3236 4920 3292
rect 4920 3236 4976 3292
rect 4976 3236 4980 3292
rect 4916 3232 4980 3236
rect 4996 3292 5060 3296
rect 4996 3236 5000 3292
rect 5000 3236 5056 3292
rect 5056 3236 5060 3292
rect 4996 3232 5060 3236
rect 5076 3292 5140 3296
rect 5076 3236 5080 3292
rect 5080 3236 5136 3292
rect 5136 3236 5140 3292
rect 5076 3232 5140 3236
rect 5156 3292 5220 3296
rect 5156 3236 5160 3292
rect 5160 3236 5216 3292
rect 5216 3236 5220 3292
rect 5156 3232 5220 3236
rect 5236 3292 5300 3296
rect 5236 3236 5240 3292
rect 5240 3236 5296 3292
rect 5296 3236 5300 3292
rect 5236 3232 5300 3236
rect 10916 3292 10980 3296
rect 10916 3236 10920 3292
rect 10920 3236 10976 3292
rect 10976 3236 10980 3292
rect 10916 3232 10980 3236
rect 10996 3292 11060 3296
rect 10996 3236 11000 3292
rect 11000 3236 11056 3292
rect 11056 3236 11060 3292
rect 10996 3232 11060 3236
rect 11076 3292 11140 3296
rect 11076 3236 11080 3292
rect 11080 3236 11136 3292
rect 11136 3236 11140 3292
rect 11076 3232 11140 3236
rect 11156 3292 11220 3296
rect 11156 3236 11160 3292
rect 11160 3236 11216 3292
rect 11216 3236 11220 3292
rect 11156 3232 11220 3236
rect 11236 3292 11300 3296
rect 11236 3236 11240 3292
rect 11240 3236 11296 3292
rect 11296 3236 11300 3292
rect 11236 3232 11300 3236
rect 16916 3292 16980 3296
rect 16916 3236 16920 3292
rect 16920 3236 16976 3292
rect 16976 3236 16980 3292
rect 16916 3232 16980 3236
rect 16996 3292 17060 3296
rect 16996 3236 17000 3292
rect 17000 3236 17056 3292
rect 17056 3236 17060 3292
rect 16996 3232 17060 3236
rect 17076 3292 17140 3296
rect 17076 3236 17080 3292
rect 17080 3236 17136 3292
rect 17136 3236 17140 3292
rect 17076 3232 17140 3236
rect 17156 3292 17220 3296
rect 17156 3236 17160 3292
rect 17160 3236 17216 3292
rect 17216 3236 17220 3292
rect 17156 3232 17220 3236
rect 17236 3292 17300 3296
rect 17236 3236 17240 3292
rect 17240 3236 17296 3292
rect 17296 3236 17300 3292
rect 17236 3232 17300 3236
rect 22916 3292 22980 3296
rect 22916 3236 22920 3292
rect 22920 3236 22976 3292
rect 22976 3236 22980 3292
rect 22916 3232 22980 3236
rect 22996 3292 23060 3296
rect 22996 3236 23000 3292
rect 23000 3236 23056 3292
rect 23056 3236 23060 3292
rect 22996 3232 23060 3236
rect 23076 3292 23140 3296
rect 23076 3236 23080 3292
rect 23080 3236 23136 3292
rect 23136 3236 23140 3292
rect 23076 3232 23140 3236
rect 23156 3292 23220 3296
rect 23156 3236 23160 3292
rect 23160 3236 23216 3292
rect 23216 3236 23220 3292
rect 23156 3232 23220 3236
rect 23236 3292 23300 3296
rect 23236 3236 23240 3292
rect 23240 3236 23296 3292
rect 23296 3236 23300 3292
rect 23236 3232 23300 3236
rect 28916 3292 28980 3296
rect 28916 3236 28920 3292
rect 28920 3236 28976 3292
rect 28976 3236 28980 3292
rect 28916 3232 28980 3236
rect 28996 3292 29060 3296
rect 28996 3236 29000 3292
rect 29000 3236 29056 3292
rect 29056 3236 29060 3292
rect 28996 3232 29060 3236
rect 29076 3292 29140 3296
rect 29076 3236 29080 3292
rect 29080 3236 29136 3292
rect 29136 3236 29140 3292
rect 29076 3232 29140 3236
rect 29156 3292 29220 3296
rect 29156 3236 29160 3292
rect 29160 3236 29216 3292
rect 29216 3236 29220 3292
rect 29156 3232 29220 3236
rect 29236 3292 29300 3296
rect 29236 3236 29240 3292
rect 29240 3236 29296 3292
rect 29296 3236 29300 3292
rect 29236 3232 29300 3236
rect 4176 2748 4240 2752
rect 4176 2692 4180 2748
rect 4180 2692 4236 2748
rect 4236 2692 4240 2748
rect 4176 2688 4240 2692
rect 4256 2748 4320 2752
rect 4256 2692 4260 2748
rect 4260 2692 4316 2748
rect 4316 2692 4320 2748
rect 4256 2688 4320 2692
rect 4336 2748 4400 2752
rect 4336 2692 4340 2748
rect 4340 2692 4396 2748
rect 4396 2692 4400 2748
rect 4336 2688 4400 2692
rect 4416 2748 4480 2752
rect 4416 2692 4420 2748
rect 4420 2692 4476 2748
rect 4476 2692 4480 2748
rect 4416 2688 4480 2692
rect 4496 2748 4560 2752
rect 4496 2692 4500 2748
rect 4500 2692 4556 2748
rect 4556 2692 4560 2748
rect 4496 2688 4560 2692
rect 10176 2748 10240 2752
rect 10176 2692 10180 2748
rect 10180 2692 10236 2748
rect 10236 2692 10240 2748
rect 10176 2688 10240 2692
rect 10256 2748 10320 2752
rect 10256 2692 10260 2748
rect 10260 2692 10316 2748
rect 10316 2692 10320 2748
rect 10256 2688 10320 2692
rect 10336 2748 10400 2752
rect 10336 2692 10340 2748
rect 10340 2692 10396 2748
rect 10396 2692 10400 2748
rect 10336 2688 10400 2692
rect 10416 2748 10480 2752
rect 10416 2692 10420 2748
rect 10420 2692 10476 2748
rect 10476 2692 10480 2748
rect 10416 2688 10480 2692
rect 10496 2748 10560 2752
rect 10496 2692 10500 2748
rect 10500 2692 10556 2748
rect 10556 2692 10560 2748
rect 10496 2688 10560 2692
rect 16176 2748 16240 2752
rect 16176 2692 16180 2748
rect 16180 2692 16236 2748
rect 16236 2692 16240 2748
rect 16176 2688 16240 2692
rect 16256 2748 16320 2752
rect 16256 2692 16260 2748
rect 16260 2692 16316 2748
rect 16316 2692 16320 2748
rect 16256 2688 16320 2692
rect 16336 2748 16400 2752
rect 16336 2692 16340 2748
rect 16340 2692 16396 2748
rect 16396 2692 16400 2748
rect 16336 2688 16400 2692
rect 16416 2748 16480 2752
rect 16416 2692 16420 2748
rect 16420 2692 16476 2748
rect 16476 2692 16480 2748
rect 16416 2688 16480 2692
rect 16496 2748 16560 2752
rect 16496 2692 16500 2748
rect 16500 2692 16556 2748
rect 16556 2692 16560 2748
rect 16496 2688 16560 2692
rect 22176 2748 22240 2752
rect 22176 2692 22180 2748
rect 22180 2692 22236 2748
rect 22236 2692 22240 2748
rect 22176 2688 22240 2692
rect 22256 2748 22320 2752
rect 22256 2692 22260 2748
rect 22260 2692 22316 2748
rect 22316 2692 22320 2748
rect 22256 2688 22320 2692
rect 22336 2748 22400 2752
rect 22336 2692 22340 2748
rect 22340 2692 22396 2748
rect 22396 2692 22400 2748
rect 22336 2688 22400 2692
rect 22416 2748 22480 2752
rect 22416 2692 22420 2748
rect 22420 2692 22476 2748
rect 22476 2692 22480 2748
rect 22416 2688 22480 2692
rect 22496 2748 22560 2752
rect 22496 2692 22500 2748
rect 22500 2692 22556 2748
rect 22556 2692 22560 2748
rect 22496 2688 22560 2692
rect 28176 2748 28240 2752
rect 28176 2692 28180 2748
rect 28180 2692 28236 2748
rect 28236 2692 28240 2748
rect 28176 2688 28240 2692
rect 28256 2748 28320 2752
rect 28256 2692 28260 2748
rect 28260 2692 28316 2748
rect 28316 2692 28320 2748
rect 28256 2688 28320 2692
rect 28336 2748 28400 2752
rect 28336 2692 28340 2748
rect 28340 2692 28396 2748
rect 28396 2692 28400 2748
rect 28336 2688 28400 2692
rect 28416 2748 28480 2752
rect 28416 2692 28420 2748
rect 28420 2692 28476 2748
rect 28476 2692 28480 2748
rect 28416 2688 28480 2692
rect 28496 2748 28560 2752
rect 28496 2692 28500 2748
rect 28500 2692 28556 2748
rect 28556 2692 28560 2748
rect 28496 2688 28560 2692
rect 14044 2484 14108 2548
rect 4916 2204 4980 2208
rect 4916 2148 4920 2204
rect 4920 2148 4976 2204
rect 4976 2148 4980 2204
rect 4916 2144 4980 2148
rect 4996 2204 5060 2208
rect 4996 2148 5000 2204
rect 5000 2148 5056 2204
rect 5056 2148 5060 2204
rect 4996 2144 5060 2148
rect 5076 2204 5140 2208
rect 5076 2148 5080 2204
rect 5080 2148 5136 2204
rect 5136 2148 5140 2204
rect 5076 2144 5140 2148
rect 5156 2204 5220 2208
rect 5156 2148 5160 2204
rect 5160 2148 5216 2204
rect 5216 2148 5220 2204
rect 5156 2144 5220 2148
rect 5236 2204 5300 2208
rect 5236 2148 5240 2204
rect 5240 2148 5296 2204
rect 5296 2148 5300 2204
rect 5236 2144 5300 2148
rect 10916 2204 10980 2208
rect 10916 2148 10920 2204
rect 10920 2148 10976 2204
rect 10976 2148 10980 2204
rect 10916 2144 10980 2148
rect 10996 2204 11060 2208
rect 10996 2148 11000 2204
rect 11000 2148 11056 2204
rect 11056 2148 11060 2204
rect 10996 2144 11060 2148
rect 11076 2204 11140 2208
rect 11076 2148 11080 2204
rect 11080 2148 11136 2204
rect 11136 2148 11140 2204
rect 11076 2144 11140 2148
rect 11156 2204 11220 2208
rect 11156 2148 11160 2204
rect 11160 2148 11216 2204
rect 11216 2148 11220 2204
rect 11156 2144 11220 2148
rect 11236 2204 11300 2208
rect 11236 2148 11240 2204
rect 11240 2148 11296 2204
rect 11296 2148 11300 2204
rect 11236 2144 11300 2148
rect 16916 2204 16980 2208
rect 16916 2148 16920 2204
rect 16920 2148 16976 2204
rect 16976 2148 16980 2204
rect 16916 2144 16980 2148
rect 16996 2204 17060 2208
rect 16996 2148 17000 2204
rect 17000 2148 17056 2204
rect 17056 2148 17060 2204
rect 16996 2144 17060 2148
rect 17076 2204 17140 2208
rect 17076 2148 17080 2204
rect 17080 2148 17136 2204
rect 17136 2148 17140 2204
rect 17076 2144 17140 2148
rect 17156 2204 17220 2208
rect 17156 2148 17160 2204
rect 17160 2148 17216 2204
rect 17216 2148 17220 2204
rect 17156 2144 17220 2148
rect 17236 2204 17300 2208
rect 17236 2148 17240 2204
rect 17240 2148 17296 2204
rect 17296 2148 17300 2204
rect 17236 2144 17300 2148
rect 22916 2204 22980 2208
rect 22916 2148 22920 2204
rect 22920 2148 22976 2204
rect 22976 2148 22980 2204
rect 22916 2144 22980 2148
rect 22996 2204 23060 2208
rect 22996 2148 23000 2204
rect 23000 2148 23056 2204
rect 23056 2148 23060 2204
rect 22996 2144 23060 2148
rect 23076 2204 23140 2208
rect 23076 2148 23080 2204
rect 23080 2148 23136 2204
rect 23136 2148 23140 2204
rect 23076 2144 23140 2148
rect 23156 2204 23220 2208
rect 23156 2148 23160 2204
rect 23160 2148 23216 2204
rect 23216 2148 23220 2204
rect 23156 2144 23220 2148
rect 23236 2204 23300 2208
rect 23236 2148 23240 2204
rect 23240 2148 23296 2204
rect 23296 2148 23300 2204
rect 23236 2144 23300 2148
rect 28916 2204 28980 2208
rect 28916 2148 28920 2204
rect 28920 2148 28976 2204
rect 28976 2148 28980 2204
rect 28916 2144 28980 2148
rect 28996 2204 29060 2208
rect 28996 2148 29000 2204
rect 29000 2148 29056 2204
rect 29056 2148 29060 2204
rect 28996 2144 29060 2148
rect 29076 2204 29140 2208
rect 29076 2148 29080 2204
rect 29080 2148 29136 2204
rect 29136 2148 29140 2204
rect 29076 2144 29140 2148
rect 29156 2204 29220 2208
rect 29156 2148 29160 2204
rect 29160 2148 29216 2204
rect 29216 2148 29220 2204
rect 29156 2144 29220 2148
rect 29236 2204 29300 2208
rect 29236 2148 29240 2204
rect 29240 2148 29296 2204
rect 29296 2148 29300 2204
rect 29236 2144 29300 2148
<< metal4 >>
rect 4168 32128 4568 32688
rect 4168 32064 4176 32128
rect 4240 32064 4256 32128
rect 4320 32064 4336 32128
rect 4400 32064 4416 32128
rect 4480 32064 4496 32128
rect 4560 32064 4568 32128
rect 4168 31040 4568 32064
rect 4168 30976 4176 31040
rect 4240 30976 4256 31040
rect 4320 30976 4336 31040
rect 4400 30976 4416 31040
rect 4480 30976 4496 31040
rect 4560 30976 4568 31040
rect 4168 29952 4568 30976
rect 4168 29888 4176 29952
rect 4240 29888 4256 29952
rect 4320 29888 4336 29952
rect 4400 29888 4416 29952
rect 4480 29888 4496 29952
rect 4560 29888 4568 29952
rect 4168 29624 4568 29888
rect 4168 29388 4250 29624
rect 4486 29388 4568 29624
rect 4168 28864 4568 29388
rect 4168 28800 4176 28864
rect 4240 28800 4256 28864
rect 4320 28800 4336 28864
rect 4400 28800 4416 28864
rect 4480 28800 4496 28864
rect 4560 28800 4568 28864
rect 4168 27776 4568 28800
rect 4168 27712 4176 27776
rect 4240 27712 4256 27776
rect 4320 27712 4336 27776
rect 4400 27712 4416 27776
rect 4480 27712 4496 27776
rect 4560 27712 4568 27776
rect 4168 26688 4568 27712
rect 4168 26624 4176 26688
rect 4240 26624 4256 26688
rect 4320 26624 4336 26688
rect 4400 26624 4416 26688
rect 4480 26624 4496 26688
rect 4560 26624 4568 26688
rect 4168 25600 4568 26624
rect 4168 25536 4176 25600
rect 4240 25536 4256 25600
rect 4320 25536 4336 25600
rect 4400 25536 4416 25600
rect 4480 25536 4496 25600
rect 4560 25536 4568 25600
rect 4168 24512 4568 25536
rect 4168 24448 4176 24512
rect 4240 24448 4256 24512
rect 4320 24448 4336 24512
rect 4400 24448 4416 24512
rect 4480 24448 4496 24512
rect 4560 24448 4568 24512
rect 4168 23624 4568 24448
rect 4168 23424 4250 23624
rect 4486 23424 4568 23624
rect 4168 23360 4176 23424
rect 4240 23388 4250 23424
rect 4486 23388 4496 23424
rect 4240 23360 4256 23388
rect 4320 23360 4336 23388
rect 4400 23360 4416 23388
rect 4480 23360 4496 23388
rect 4560 23360 4568 23424
rect 4168 22336 4568 23360
rect 4168 22272 4176 22336
rect 4240 22272 4256 22336
rect 4320 22272 4336 22336
rect 4400 22272 4416 22336
rect 4480 22272 4496 22336
rect 4560 22272 4568 22336
rect 4168 21248 4568 22272
rect 4168 21184 4176 21248
rect 4240 21184 4256 21248
rect 4320 21184 4336 21248
rect 4400 21184 4416 21248
rect 4480 21184 4496 21248
rect 4560 21184 4568 21248
rect 4168 20160 4568 21184
rect 4168 20096 4176 20160
rect 4240 20096 4256 20160
rect 4320 20096 4336 20160
rect 4400 20096 4416 20160
rect 4480 20096 4496 20160
rect 4560 20096 4568 20160
rect 4168 19072 4568 20096
rect 4168 19008 4176 19072
rect 4240 19008 4256 19072
rect 4320 19008 4336 19072
rect 4400 19008 4416 19072
rect 4480 19008 4496 19072
rect 4560 19008 4568 19072
rect 4168 17984 4568 19008
rect 4168 17920 4176 17984
rect 4240 17920 4256 17984
rect 4320 17920 4336 17984
rect 4400 17920 4416 17984
rect 4480 17920 4496 17984
rect 4560 17920 4568 17984
rect 4168 17624 4568 17920
rect 4168 17388 4250 17624
rect 4486 17388 4568 17624
rect 4168 16896 4568 17388
rect 4168 16832 4176 16896
rect 4240 16832 4256 16896
rect 4320 16832 4336 16896
rect 4400 16832 4416 16896
rect 4480 16832 4496 16896
rect 4560 16832 4568 16896
rect 4168 15808 4568 16832
rect 4168 15744 4176 15808
rect 4240 15744 4256 15808
rect 4320 15744 4336 15808
rect 4400 15744 4416 15808
rect 4480 15744 4496 15808
rect 4560 15744 4568 15808
rect 4168 14720 4568 15744
rect 4168 14656 4176 14720
rect 4240 14656 4256 14720
rect 4320 14656 4336 14720
rect 4400 14656 4416 14720
rect 4480 14656 4496 14720
rect 4560 14656 4568 14720
rect 4168 13632 4568 14656
rect 4168 13568 4176 13632
rect 4240 13568 4256 13632
rect 4320 13568 4336 13632
rect 4400 13568 4416 13632
rect 4480 13568 4496 13632
rect 4560 13568 4568 13632
rect 4168 12544 4568 13568
rect 4168 12480 4176 12544
rect 4240 12480 4256 12544
rect 4320 12480 4336 12544
rect 4400 12480 4416 12544
rect 4480 12480 4496 12544
rect 4560 12480 4568 12544
rect 4168 11624 4568 12480
rect 4168 11456 4250 11624
rect 4486 11456 4568 11624
rect 4168 11392 4176 11456
rect 4240 11392 4250 11456
rect 4486 11392 4496 11456
rect 4560 11392 4568 11456
rect 4168 11388 4250 11392
rect 4486 11388 4568 11392
rect 4168 10368 4568 11388
rect 4168 10304 4176 10368
rect 4240 10304 4256 10368
rect 4320 10304 4336 10368
rect 4400 10304 4416 10368
rect 4480 10304 4496 10368
rect 4560 10304 4568 10368
rect 4168 9280 4568 10304
rect 4168 9216 4176 9280
rect 4240 9216 4256 9280
rect 4320 9216 4336 9280
rect 4400 9216 4416 9280
rect 4480 9216 4496 9280
rect 4560 9216 4568 9280
rect 4168 8192 4568 9216
rect 4168 8128 4176 8192
rect 4240 8128 4256 8192
rect 4320 8128 4336 8192
rect 4400 8128 4416 8192
rect 4480 8128 4496 8192
rect 4560 8128 4568 8192
rect 4168 7104 4568 8128
rect 4168 7040 4176 7104
rect 4240 7040 4256 7104
rect 4320 7040 4336 7104
rect 4400 7040 4416 7104
rect 4480 7040 4496 7104
rect 4560 7040 4568 7104
rect 4168 6016 4568 7040
rect 4168 5952 4176 6016
rect 4240 5952 4256 6016
rect 4320 5952 4336 6016
rect 4400 5952 4416 6016
rect 4480 5952 4496 6016
rect 4560 5952 4568 6016
rect 4168 5624 4568 5952
rect 4168 5388 4250 5624
rect 4486 5388 4568 5624
rect 4168 4928 4568 5388
rect 4168 4864 4176 4928
rect 4240 4864 4256 4928
rect 4320 4864 4336 4928
rect 4400 4864 4416 4928
rect 4480 4864 4496 4928
rect 4560 4864 4568 4928
rect 4168 3840 4568 4864
rect 4168 3776 4176 3840
rect 4240 3776 4256 3840
rect 4320 3776 4336 3840
rect 4400 3776 4416 3840
rect 4480 3776 4496 3840
rect 4560 3776 4568 3840
rect 4168 2752 4568 3776
rect 4168 2688 4176 2752
rect 4240 2688 4256 2752
rect 4320 2688 4336 2752
rect 4400 2688 4416 2752
rect 4480 2688 4496 2752
rect 4560 2688 4568 2752
rect 4168 2128 4568 2688
rect 4908 32672 5308 32688
rect 4908 32608 4916 32672
rect 4980 32608 4996 32672
rect 5060 32608 5076 32672
rect 5140 32608 5156 32672
rect 5220 32608 5236 32672
rect 5300 32608 5308 32672
rect 4908 31584 5308 32608
rect 4908 31520 4916 31584
rect 4980 31520 4996 31584
rect 5060 31520 5076 31584
rect 5140 31520 5156 31584
rect 5220 31520 5236 31584
rect 5300 31520 5308 31584
rect 4908 30496 5308 31520
rect 4908 30432 4916 30496
rect 4980 30432 4996 30496
rect 5060 30432 5076 30496
rect 5140 30432 5156 30496
rect 5220 30432 5236 30496
rect 5300 30432 5308 30496
rect 4908 30364 5308 30432
rect 4908 30128 4990 30364
rect 5226 30128 5308 30364
rect 4908 29408 5308 30128
rect 4908 29344 4916 29408
rect 4980 29344 4996 29408
rect 5060 29344 5076 29408
rect 5140 29344 5156 29408
rect 5220 29344 5236 29408
rect 5300 29344 5308 29408
rect 4908 28320 5308 29344
rect 4908 28256 4916 28320
rect 4980 28256 4996 28320
rect 5060 28256 5076 28320
rect 5140 28256 5156 28320
rect 5220 28256 5236 28320
rect 5300 28256 5308 28320
rect 4908 27232 5308 28256
rect 4908 27168 4916 27232
rect 4980 27168 4996 27232
rect 5060 27168 5076 27232
rect 5140 27168 5156 27232
rect 5220 27168 5236 27232
rect 5300 27168 5308 27232
rect 4908 26144 5308 27168
rect 4908 26080 4916 26144
rect 4980 26080 4996 26144
rect 5060 26080 5076 26144
rect 5140 26080 5156 26144
rect 5220 26080 5236 26144
rect 5300 26080 5308 26144
rect 4908 25056 5308 26080
rect 4908 24992 4916 25056
rect 4980 24992 4996 25056
rect 5060 24992 5076 25056
rect 5140 24992 5156 25056
rect 5220 24992 5236 25056
rect 5300 24992 5308 25056
rect 4908 24364 5308 24992
rect 4908 24128 4990 24364
rect 5226 24128 5308 24364
rect 4908 23968 5308 24128
rect 4908 23904 4916 23968
rect 4980 23904 4996 23968
rect 5060 23904 5076 23968
rect 5140 23904 5156 23968
rect 5220 23904 5236 23968
rect 5300 23904 5308 23968
rect 4908 22880 5308 23904
rect 4908 22816 4916 22880
rect 4980 22816 4996 22880
rect 5060 22816 5076 22880
rect 5140 22816 5156 22880
rect 5220 22816 5236 22880
rect 5300 22816 5308 22880
rect 4908 21792 5308 22816
rect 4908 21728 4916 21792
rect 4980 21728 4996 21792
rect 5060 21728 5076 21792
rect 5140 21728 5156 21792
rect 5220 21728 5236 21792
rect 5300 21728 5308 21792
rect 4908 20704 5308 21728
rect 4908 20640 4916 20704
rect 4980 20640 4996 20704
rect 5060 20640 5076 20704
rect 5140 20640 5156 20704
rect 5220 20640 5236 20704
rect 5300 20640 5308 20704
rect 4908 19616 5308 20640
rect 4908 19552 4916 19616
rect 4980 19552 4996 19616
rect 5060 19552 5076 19616
rect 5140 19552 5156 19616
rect 5220 19552 5236 19616
rect 5300 19552 5308 19616
rect 4908 18528 5308 19552
rect 4908 18464 4916 18528
rect 4980 18464 4996 18528
rect 5060 18464 5076 18528
rect 5140 18464 5156 18528
rect 5220 18464 5236 18528
rect 5300 18464 5308 18528
rect 4908 18364 5308 18464
rect 4908 18128 4990 18364
rect 5226 18128 5308 18364
rect 4908 17440 5308 18128
rect 4908 17376 4916 17440
rect 4980 17376 4996 17440
rect 5060 17376 5076 17440
rect 5140 17376 5156 17440
rect 5220 17376 5236 17440
rect 5300 17376 5308 17440
rect 4908 16352 5308 17376
rect 4908 16288 4916 16352
rect 4980 16288 4996 16352
rect 5060 16288 5076 16352
rect 5140 16288 5156 16352
rect 5220 16288 5236 16352
rect 5300 16288 5308 16352
rect 4908 15264 5308 16288
rect 4908 15200 4916 15264
rect 4980 15200 4996 15264
rect 5060 15200 5076 15264
rect 5140 15200 5156 15264
rect 5220 15200 5236 15264
rect 5300 15200 5308 15264
rect 4908 14176 5308 15200
rect 4908 14112 4916 14176
rect 4980 14112 4996 14176
rect 5060 14112 5076 14176
rect 5140 14112 5156 14176
rect 5220 14112 5236 14176
rect 5300 14112 5308 14176
rect 4908 13088 5308 14112
rect 4908 13024 4916 13088
rect 4980 13024 4996 13088
rect 5060 13024 5076 13088
rect 5140 13024 5156 13088
rect 5220 13024 5236 13088
rect 5300 13024 5308 13088
rect 4908 12364 5308 13024
rect 4908 12128 4990 12364
rect 5226 12128 5308 12364
rect 4908 12000 5308 12128
rect 4908 11936 4916 12000
rect 4980 11936 4996 12000
rect 5060 11936 5076 12000
rect 5140 11936 5156 12000
rect 5220 11936 5236 12000
rect 5300 11936 5308 12000
rect 4908 10912 5308 11936
rect 4908 10848 4916 10912
rect 4980 10848 4996 10912
rect 5060 10848 5076 10912
rect 5140 10848 5156 10912
rect 5220 10848 5236 10912
rect 5300 10848 5308 10912
rect 4908 9824 5308 10848
rect 4908 9760 4916 9824
rect 4980 9760 4996 9824
rect 5060 9760 5076 9824
rect 5140 9760 5156 9824
rect 5220 9760 5236 9824
rect 5300 9760 5308 9824
rect 4908 8736 5308 9760
rect 4908 8672 4916 8736
rect 4980 8672 4996 8736
rect 5060 8672 5076 8736
rect 5140 8672 5156 8736
rect 5220 8672 5236 8736
rect 5300 8672 5308 8736
rect 4908 7648 5308 8672
rect 10168 32128 10568 32688
rect 10168 32064 10176 32128
rect 10240 32064 10256 32128
rect 10320 32064 10336 32128
rect 10400 32064 10416 32128
rect 10480 32064 10496 32128
rect 10560 32064 10568 32128
rect 10168 31040 10568 32064
rect 10168 30976 10176 31040
rect 10240 30976 10256 31040
rect 10320 30976 10336 31040
rect 10400 30976 10416 31040
rect 10480 30976 10496 31040
rect 10560 30976 10568 31040
rect 10168 29952 10568 30976
rect 10168 29888 10176 29952
rect 10240 29888 10256 29952
rect 10320 29888 10336 29952
rect 10400 29888 10416 29952
rect 10480 29888 10496 29952
rect 10560 29888 10568 29952
rect 10168 29624 10568 29888
rect 10168 29388 10250 29624
rect 10486 29388 10568 29624
rect 10168 28864 10568 29388
rect 10168 28800 10176 28864
rect 10240 28800 10256 28864
rect 10320 28800 10336 28864
rect 10400 28800 10416 28864
rect 10480 28800 10496 28864
rect 10560 28800 10568 28864
rect 10168 27776 10568 28800
rect 10168 27712 10176 27776
rect 10240 27712 10256 27776
rect 10320 27712 10336 27776
rect 10400 27712 10416 27776
rect 10480 27712 10496 27776
rect 10560 27712 10568 27776
rect 10168 26688 10568 27712
rect 10168 26624 10176 26688
rect 10240 26624 10256 26688
rect 10320 26624 10336 26688
rect 10400 26624 10416 26688
rect 10480 26624 10496 26688
rect 10560 26624 10568 26688
rect 10168 25600 10568 26624
rect 10168 25536 10176 25600
rect 10240 25536 10256 25600
rect 10320 25536 10336 25600
rect 10400 25536 10416 25600
rect 10480 25536 10496 25600
rect 10560 25536 10568 25600
rect 10168 24512 10568 25536
rect 10168 24448 10176 24512
rect 10240 24448 10256 24512
rect 10320 24448 10336 24512
rect 10400 24448 10416 24512
rect 10480 24448 10496 24512
rect 10560 24448 10568 24512
rect 10168 23624 10568 24448
rect 10168 23424 10250 23624
rect 10486 23424 10568 23624
rect 10168 23360 10176 23424
rect 10240 23388 10250 23424
rect 10486 23388 10496 23424
rect 10240 23360 10256 23388
rect 10320 23360 10336 23388
rect 10400 23360 10416 23388
rect 10480 23360 10496 23388
rect 10560 23360 10568 23424
rect 10168 22336 10568 23360
rect 10168 22272 10176 22336
rect 10240 22272 10256 22336
rect 10320 22272 10336 22336
rect 10400 22272 10416 22336
rect 10480 22272 10496 22336
rect 10560 22272 10568 22336
rect 10168 21248 10568 22272
rect 10168 21184 10176 21248
rect 10240 21184 10256 21248
rect 10320 21184 10336 21248
rect 10400 21184 10416 21248
rect 10480 21184 10496 21248
rect 10560 21184 10568 21248
rect 10168 20160 10568 21184
rect 10168 20096 10176 20160
rect 10240 20096 10256 20160
rect 10320 20096 10336 20160
rect 10400 20096 10416 20160
rect 10480 20096 10496 20160
rect 10560 20096 10568 20160
rect 10168 19072 10568 20096
rect 10168 19008 10176 19072
rect 10240 19008 10256 19072
rect 10320 19008 10336 19072
rect 10400 19008 10416 19072
rect 10480 19008 10496 19072
rect 10560 19008 10568 19072
rect 10168 17984 10568 19008
rect 10168 17920 10176 17984
rect 10240 17920 10256 17984
rect 10320 17920 10336 17984
rect 10400 17920 10416 17984
rect 10480 17920 10496 17984
rect 10560 17920 10568 17984
rect 10168 17624 10568 17920
rect 10168 17388 10250 17624
rect 10486 17388 10568 17624
rect 10168 16896 10568 17388
rect 10168 16832 10176 16896
rect 10240 16832 10256 16896
rect 10320 16832 10336 16896
rect 10400 16832 10416 16896
rect 10480 16832 10496 16896
rect 10560 16832 10568 16896
rect 10168 15808 10568 16832
rect 10168 15744 10176 15808
rect 10240 15744 10256 15808
rect 10320 15744 10336 15808
rect 10400 15744 10416 15808
rect 10480 15744 10496 15808
rect 10560 15744 10568 15808
rect 10168 14720 10568 15744
rect 10168 14656 10176 14720
rect 10240 14656 10256 14720
rect 10320 14656 10336 14720
rect 10400 14656 10416 14720
rect 10480 14656 10496 14720
rect 10560 14656 10568 14720
rect 10168 13632 10568 14656
rect 10168 13568 10176 13632
rect 10240 13568 10256 13632
rect 10320 13568 10336 13632
rect 10400 13568 10416 13632
rect 10480 13568 10496 13632
rect 10560 13568 10568 13632
rect 10168 12544 10568 13568
rect 10168 12480 10176 12544
rect 10240 12480 10256 12544
rect 10320 12480 10336 12544
rect 10400 12480 10416 12544
rect 10480 12480 10496 12544
rect 10560 12480 10568 12544
rect 10168 11624 10568 12480
rect 10168 11456 10250 11624
rect 10486 11456 10568 11624
rect 10168 11392 10176 11456
rect 10240 11392 10250 11456
rect 10486 11392 10496 11456
rect 10560 11392 10568 11456
rect 10168 11388 10250 11392
rect 10486 11388 10568 11392
rect 10168 10368 10568 11388
rect 10168 10304 10176 10368
rect 10240 10304 10256 10368
rect 10320 10304 10336 10368
rect 10400 10304 10416 10368
rect 10480 10304 10496 10368
rect 10560 10304 10568 10368
rect 10168 9280 10568 10304
rect 10168 9216 10176 9280
rect 10240 9216 10256 9280
rect 10320 9216 10336 9280
rect 10400 9216 10416 9280
rect 10480 9216 10496 9280
rect 10560 9216 10568 9280
rect 9995 8532 10061 8533
rect 9995 8468 9996 8532
rect 10060 8468 10061 8532
rect 9995 8467 10061 8468
rect 4908 7584 4916 7648
rect 4980 7584 4996 7648
rect 5060 7584 5076 7648
rect 5140 7584 5156 7648
rect 5220 7584 5236 7648
rect 5300 7584 5308 7648
rect 4908 6560 5308 7584
rect 4908 6496 4916 6560
rect 4980 6496 4996 6560
rect 5060 6496 5076 6560
rect 5140 6496 5156 6560
rect 5220 6496 5236 6560
rect 5300 6496 5308 6560
rect 4908 6364 5308 6496
rect 4908 6128 4990 6364
rect 5226 6128 5308 6364
rect 4908 5472 5308 6128
rect 4908 5408 4916 5472
rect 4980 5408 4996 5472
rect 5060 5408 5076 5472
rect 5140 5408 5156 5472
rect 5220 5408 5236 5472
rect 5300 5408 5308 5472
rect 4908 4384 5308 5408
rect 9998 4997 10058 8467
rect 10168 8192 10568 9216
rect 10908 32672 11308 32688
rect 10908 32608 10916 32672
rect 10980 32608 10996 32672
rect 11060 32608 11076 32672
rect 11140 32608 11156 32672
rect 11220 32608 11236 32672
rect 11300 32608 11308 32672
rect 10908 31584 11308 32608
rect 10908 31520 10916 31584
rect 10980 31520 10996 31584
rect 11060 31520 11076 31584
rect 11140 31520 11156 31584
rect 11220 31520 11236 31584
rect 11300 31520 11308 31584
rect 10908 30496 11308 31520
rect 10908 30432 10916 30496
rect 10980 30432 10996 30496
rect 11060 30432 11076 30496
rect 11140 30432 11156 30496
rect 11220 30432 11236 30496
rect 11300 30432 11308 30496
rect 10908 30364 11308 30432
rect 10908 30128 10990 30364
rect 11226 30128 11308 30364
rect 10908 29408 11308 30128
rect 10908 29344 10916 29408
rect 10980 29344 10996 29408
rect 11060 29344 11076 29408
rect 11140 29344 11156 29408
rect 11220 29344 11236 29408
rect 11300 29344 11308 29408
rect 10908 28320 11308 29344
rect 16168 32128 16568 32688
rect 16168 32064 16176 32128
rect 16240 32064 16256 32128
rect 16320 32064 16336 32128
rect 16400 32064 16416 32128
rect 16480 32064 16496 32128
rect 16560 32064 16568 32128
rect 16168 31040 16568 32064
rect 16168 30976 16176 31040
rect 16240 30976 16256 31040
rect 16320 30976 16336 31040
rect 16400 30976 16416 31040
rect 16480 30976 16496 31040
rect 16560 30976 16568 31040
rect 16168 29952 16568 30976
rect 16168 29888 16176 29952
rect 16240 29888 16256 29952
rect 16320 29888 16336 29952
rect 16400 29888 16416 29952
rect 16480 29888 16496 29952
rect 16560 29888 16568 29952
rect 16168 29624 16568 29888
rect 16168 29388 16250 29624
rect 16486 29388 16568 29624
rect 14043 29068 14109 29069
rect 14043 29004 14044 29068
rect 14108 29004 14109 29068
rect 14043 29003 14109 29004
rect 10908 28256 10916 28320
rect 10980 28256 10996 28320
rect 11060 28256 11076 28320
rect 11140 28256 11156 28320
rect 11220 28256 11236 28320
rect 11300 28256 11308 28320
rect 10908 27232 11308 28256
rect 10908 27168 10916 27232
rect 10980 27168 10996 27232
rect 11060 27168 11076 27232
rect 11140 27168 11156 27232
rect 11220 27168 11236 27232
rect 11300 27168 11308 27232
rect 10908 26144 11308 27168
rect 10908 26080 10916 26144
rect 10980 26080 10996 26144
rect 11060 26080 11076 26144
rect 11140 26080 11156 26144
rect 11220 26080 11236 26144
rect 11300 26080 11308 26144
rect 10908 25056 11308 26080
rect 10908 24992 10916 25056
rect 10980 24992 10996 25056
rect 11060 24992 11076 25056
rect 11140 24992 11156 25056
rect 11220 24992 11236 25056
rect 11300 24992 11308 25056
rect 10908 24364 11308 24992
rect 10908 24128 10990 24364
rect 11226 24128 11308 24364
rect 10908 23968 11308 24128
rect 10908 23904 10916 23968
rect 10980 23904 10996 23968
rect 11060 23904 11076 23968
rect 11140 23904 11156 23968
rect 11220 23904 11236 23968
rect 11300 23904 11308 23968
rect 10908 22880 11308 23904
rect 10908 22816 10916 22880
rect 10980 22816 10996 22880
rect 11060 22816 11076 22880
rect 11140 22816 11156 22880
rect 11220 22816 11236 22880
rect 11300 22816 11308 22880
rect 10908 21792 11308 22816
rect 10908 21728 10916 21792
rect 10980 21728 10996 21792
rect 11060 21728 11076 21792
rect 11140 21728 11156 21792
rect 11220 21728 11236 21792
rect 11300 21728 11308 21792
rect 10908 20704 11308 21728
rect 12939 20772 13005 20773
rect 12939 20708 12940 20772
rect 13004 20708 13005 20772
rect 12939 20707 13005 20708
rect 10908 20640 10916 20704
rect 10980 20640 10996 20704
rect 11060 20640 11076 20704
rect 11140 20640 11156 20704
rect 11220 20640 11236 20704
rect 11300 20640 11308 20704
rect 10908 19616 11308 20640
rect 10908 19552 10916 19616
rect 10980 19552 10996 19616
rect 11060 19552 11076 19616
rect 11140 19552 11156 19616
rect 11220 19552 11236 19616
rect 11300 19552 11308 19616
rect 10908 18528 11308 19552
rect 10908 18464 10916 18528
rect 10980 18464 10996 18528
rect 11060 18464 11076 18528
rect 11140 18464 11156 18528
rect 11220 18464 11236 18528
rect 11300 18464 11308 18528
rect 10908 18364 11308 18464
rect 10908 18128 10990 18364
rect 11226 18128 11308 18364
rect 10908 17440 11308 18128
rect 10908 17376 10916 17440
rect 10980 17376 10996 17440
rect 11060 17376 11076 17440
rect 11140 17376 11156 17440
rect 11220 17376 11236 17440
rect 11300 17376 11308 17440
rect 10908 16352 11308 17376
rect 10908 16288 10916 16352
rect 10980 16288 10996 16352
rect 11060 16288 11076 16352
rect 11140 16288 11156 16352
rect 11220 16288 11236 16352
rect 11300 16288 11308 16352
rect 10908 15264 11308 16288
rect 10908 15200 10916 15264
rect 10980 15200 10996 15264
rect 11060 15200 11076 15264
rect 11140 15200 11156 15264
rect 11220 15200 11236 15264
rect 11300 15200 11308 15264
rect 10908 14176 11308 15200
rect 10908 14112 10916 14176
rect 10980 14112 10996 14176
rect 11060 14112 11076 14176
rect 11140 14112 11156 14176
rect 11220 14112 11236 14176
rect 11300 14112 11308 14176
rect 10908 13088 11308 14112
rect 10908 13024 10916 13088
rect 10980 13024 10996 13088
rect 11060 13024 11076 13088
rect 11140 13024 11156 13088
rect 11220 13024 11236 13088
rect 11300 13024 11308 13088
rect 10908 12364 11308 13024
rect 12942 12749 13002 20707
rect 12939 12748 13005 12749
rect 12939 12684 12940 12748
rect 13004 12684 13005 12748
rect 12939 12683 13005 12684
rect 10908 12128 10990 12364
rect 11226 12128 11308 12364
rect 10908 12000 11308 12128
rect 10908 11936 10916 12000
rect 10980 11936 10996 12000
rect 11060 11936 11076 12000
rect 11140 11936 11156 12000
rect 11220 11936 11236 12000
rect 11300 11936 11308 12000
rect 10908 10912 11308 11936
rect 12942 11389 13002 12683
rect 12939 11388 13005 11389
rect 12939 11324 12940 11388
rect 13004 11324 13005 11388
rect 12939 11323 13005 11324
rect 10908 10848 10916 10912
rect 10980 10848 10996 10912
rect 11060 10848 11076 10912
rect 11140 10848 11156 10912
rect 11220 10848 11236 10912
rect 11300 10848 11308 10912
rect 10908 9824 11308 10848
rect 10908 9760 10916 9824
rect 10980 9760 10996 9824
rect 11060 9760 11076 9824
rect 11140 9760 11156 9824
rect 11220 9760 11236 9824
rect 11300 9760 11308 9824
rect 10731 8940 10797 8941
rect 10731 8876 10732 8940
rect 10796 8876 10797 8940
rect 10731 8875 10797 8876
rect 10168 8128 10176 8192
rect 10240 8128 10256 8192
rect 10320 8128 10336 8192
rect 10400 8128 10416 8192
rect 10480 8128 10496 8192
rect 10560 8128 10568 8192
rect 10168 7104 10568 8128
rect 10168 7040 10176 7104
rect 10240 7040 10256 7104
rect 10320 7040 10336 7104
rect 10400 7040 10416 7104
rect 10480 7040 10496 7104
rect 10560 7040 10568 7104
rect 10168 6016 10568 7040
rect 10734 6765 10794 8875
rect 10908 8736 11308 9760
rect 10908 8672 10916 8736
rect 10980 8672 10996 8736
rect 11060 8672 11076 8736
rect 11140 8672 11156 8736
rect 11220 8672 11236 8736
rect 11300 8672 11308 8736
rect 10908 7648 11308 8672
rect 10908 7584 10916 7648
rect 10980 7584 10996 7648
rect 11060 7584 11076 7648
rect 11140 7584 11156 7648
rect 11220 7584 11236 7648
rect 11300 7584 11308 7648
rect 10731 6764 10797 6765
rect 10731 6700 10732 6764
rect 10796 6700 10797 6764
rect 10731 6699 10797 6700
rect 10168 5952 10176 6016
rect 10240 5952 10256 6016
rect 10320 5952 10336 6016
rect 10400 5952 10416 6016
rect 10480 5952 10496 6016
rect 10560 5952 10568 6016
rect 10168 5624 10568 5952
rect 10168 5388 10250 5624
rect 10486 5388 10568 5624
rect 9995 4996 10061 4997
rect 9995 4932 9996 4996
rect 10060 4932 10061 4996
rect 9995 4931 10061 4932
rect 4908 4320 4916 4384
rect 4980 4320 4996 4384
rect 5060 4320 5076 4384
rect 5140 4320 5156 4384
rect 5220 4320 5236 4384
rect 5300 4320 5308 4384
rect 4908 3296 5308 4320
rect 4908 3232 4916 3296
rect 4980 3232 4996 3296
rect 5060 3232 5076 3296
rect 5140 3232 5156 3296
rect 5220 3232 5236 3296
rect 5300 3232 5308 3296
rect 4908 2208 5308 3232
rect 4908 2144 4916 2208
rect 4980 2144 4996 2208
rect 5060 2144 5076 2208
rect 5140 2144 5156 2208
rect 5220 2144 5236 2208
rect 5300 2144 5308 2208
rect 4908 2128 5308 2144
rect 10168 4928 10568 5388
rect 10168 4864 10176 4928
rect 10240 4864 10256 4928
rect 10320 4864 10336 4928
rect 10400 4864 10416 4928
rect 10480 4864 10496 4928
rect 10560 4864 10568 4928
rect 10168 3840 10568 4864
rect 10168 3776 10176 3840
rect 10240 3776 10256 3840
rect 10320 3776 10336 3840
rect 10400 3776 10416 3840
rect 10480 3776 10496 3840
rect 10560 3776 10568 3840
rect 10168 2752 10568 3776
rect 10168 2688 10176 2752
rect 10240 2688 10256 2752
rect 10320 2688 10336 2752
rect 10400 2688 10416 2752
rect 10480 2688 10496 2752
rect 10560 2688 10568 2752
rect 10168 2128 10568 2688
rect 10908 6560 11308 7584
rect 10908 6496 10916 6560
rect 10980 6496 10996 6560
rect 11060 6496 11076 6560
rect 11140 6496 11156 6560
rect 11220 6496 11236 6560
rect 11300 6496 11308 6560
rect 10908 6364 11308 6496
rect 10908 6128 10990 6364
rect 11226 6128 11308 6364
rect 10908 5472 11308 6128
rect 10908 5408 10916 5472
rect 10980 5408 10996 5472
rect 11060 5408 11076 5472
rect 11140 5408 11156 5472
rect 11220 5408 11236 5472
rect 11300 5408 11308 5472
rect 10908 4384 11308 5408
rect 10908 4320 10916 4384
rect 10980 4320 10996 4384
rect 11060 4320 11076 4384
rect 11140 4320 11156 4384
rect 11220 4320 11236 4384
rect 11300 4320 11308 4384
rect 10908 3296 11308 4320
rect 10908 3232 10916 3296
rect 10980 3232 10996 3296
rect 11060 3232 11076 3296
rect 11140 3232 11156 3296
rect 11220 3232 11236 3296
rect 11300 3232 11308 3296
rect 10908 2208 11308 3232
rect 14046 2549 14106 29003
rect 16168 28864 16568 29388
rect 16168 28800 16176 28864
rect 16240 28800 16256 28864
rect 16320 28800 16336 28864
rect 16400 28800 16416 28864
rect 16480 28800 16496 28864
rect 16560 28800 16568 28864
rect 16168 27776 16568 28800
rect 16168 27712 16176 27776
rect 16240 27712 16256 27776
rect 16320 27712 16336 27776
rect 16400 27712 16416 27776
rect 16480 27712 16496 27776
rect 16560 27712 16568 27776
rect 16168 26688 16568 27712
rect 16168 26624 16176 26688
rect 16240 26624 16256 26688
rect 16320 26624 16336 26688
rect 16400 26624 16416 26688
rect 16480 26624 16496 26688
rect 16560 26624 16568 26688
rect 16168 25600 16568 26624
rect 16168 25536 16176 25600
rect 16240 25536 16256 25600
rect 16320 25536 16336 25600
rect 16400 25536 16416 25600
rect 16480 25536 16496 25600
rect 16560 25536 16568 25600
rect 16168 24512 16568 25536
rect 16168 24448 16176 24512
rect 16240 24448 16256 24512
rect 16320 24448 16336 24512
rect 16400 24448 16416 24512
rect 16480 24448 16496 24512
rect 16560 24448 16568 24512
rect 16168 23624 16568 24448
rect 14227 23492 14293 23493
rect 14227 23428 14228 23492
rect 14292 23428 14293 23492
rect 14227 23427 14293 23428
rect 14230 19413 14290 23427
rect 16168 23424 16250 23624
rect 16486 23424 16568 23624
rect 16168 23360 16176 23424
rect 16240 23388 16250 23424
rect 16486 23388 16496 23424
rect 16240 23360 16256 23388
rect 16320 23360 16336 23388
rect 16400 23360 16416 23388
rect 16480 23360 16496 23388
rect 16560 23360 16568 23424
rect 16168 22336 16568 23360
rect 16168 22272 16176 22336
rect 16240 22272 16256 22336
rect 16320 22272 16336 22336
rect 16400 22272 16416 22336
rect 16480 22272 16496 22336
rect 16560 22272 16568 22336
rect 16168 21248 16568 22272
rect 16168 21184 16176 21248
rect 16240 21184 16256 21248
rect 16320 21184 16336 21248
rect 16400 21184 16416 21248
rect 16480 21184 16496 21248
rect 16560 21184 16568 21248
rect 16168 20160 16568 21184
rect 16168 20096 16176 20160
rect 16240 20096 16256 20160
rect 16320 20096 16336 20160
rect 16400 20096 16416 20160
rect 16480 20096 16496 20160
rect 16560 20096 16568 20160
rect 14227 19412 14293 19413
rect 14227 19348 14228 19412
rect 14292 19348 14293 19412
rect 14227 19347 14293 19348
rect 16168 19072 16568 20096
rect 16168 19008 16176 19072
rect 16240 19008 16256 19072
rect 16320 19008 16336 19072
rect 16400 19008 16416 19072
rect 16480 19008 16496 19072
rect 16560 19008 16568 19072
rect 16168 17984 16568 19008
rect 16168 17920 16176 17984
rect 16240 17920 16256 17984
rect 16320 17920 16336 17984
rect 16400 17920 16416 17984
rect 16480 17920 16496 17984
rect 16560 17920 16568 17984
rect 16168 17624 16568 17920
rect 16168 17388 16250 17624
rect 16486 17388 16568 17624
rect 16168 16896 16568 17388
rect 16168 16832 16176 16896
rect 16240 16832 16256 16896
rect 16320 16832 16336 16896
rect 16400 16832 16416 16896
rect 16480 16832 16496 16896
rect 16560 16832 16568 16896
rect 16168 15808 16568 16832
rect 16168 15744 16176 15808
rect 16240 15744 16256 15808
rect 16320 15744 16336 15808
rect 16400 15744 16416 15808
rect 16480 15744 16496 15808
rect 16560 15744 16568 15808
rect 16168 14720 16568 15744
rect 16168 14656 16176 14720
rect 16240 14656 16256 14720
rect 16320 14656 16336 14720
rect 16400 14656 16416 14720
rect 16480 14656 16496 14720
rect 16560 14656 16568 14720
rect 16168 13632 16568 14656
rect 16168 13568 16176 13632
rect 16240 13568 16256 13632
rect 16320 13568 16336 13632
rect 16400 13568 16416 13632
rect 16480 13568 16496 13632
rect 16560 13568 16568 13632
rect 16168 12544 16568 13568
rect 16168 12480 16176 12544
rect 16240 12480 16256 12544
rect 16320 12480 16336 12544
rect 16400 12480 16416 12544
rect 16480 12480 16496 12544
rect 16560 12480 16568 12544
rect 16168 11624 16568 12480
rect 16168 11456 16250 11624
rect 16486 11456 16568 11624
rect 16168 11392 16176 11456
rect 16240 11392 16250 11456
rect 16486 11392 16496 11456
rect 16560 11392 16568 11456
rect 16168 11388 16250 11392
rect 16486 11388 16568 11392
rect 16168 10368 16568 11388
rect 16168 10304 16176 10368
rect 16240 10304 16256 10368
rect 16320 10304 16336 10368
rect 16400 10304 16416 10368
rect 16480 10304 16496 10368
rect 16560 10304 16568 10368
rect 16168 9280 16568 10304
rect 16168 9216 16176 9280
rect 16240 9216 16256 9280
rect 16320 9216 16336 9280
rect 16400 9216 16416 9280
rect 16480 9216 16496 9280
rect 16560 9216 16568 9280
rect 16168 8192 16568 9216
rect 16168 8128 16176 8192
rect 16240 8128 16256 8192
rect 16320 8128 16336 8192
rect 16400 8128 16416 8192
rect 16480 8128 16496 8192
rect 16560 8128 16568 8192
rect 16168 7104 16568 8128
rect 16168 7040 16176 7104
rect 16240 7040 16256 7104
rect 16320 7040 16336 7104
rect 16400 7040 16416 7104
rect 16480 7040 16496 7104
rect 16560 7040 16568 7104
rect 16168 6016 16568 7040
rect 16168 5952 16176 6016
rect 16240 5952 16256 6016
rect 16320 5952 16336 6016
rect 16400 5952 16416 6016
rect 16480 5952 16496 6016
rect 16560 5952 16568 6016
rect 16168 5624 16568 5952
rect 16168 5388 16250 5624
rect 16486 5388 16568 5624
rect 16168 4928 16568 5388
rect 16168 4864 16176 4928
rect 16240 4864 16256 4928
rect 16320 4864 16336 4928
rect 16400 4864 16416 4928
rect 16480 4864 16496 4928
rect 16560 4864 16568 4928
rect 16168 3840 16568 4864
rect 16168 3776 16176 3840
rect 16240 3776 16256 3840
rect 16320 3776 16336 3840
rect 16400 3776 16416 3840
rect 16480 3776 16496 3840
rect 16560 3776 16568 3840
rect 16168 2752 16568 3776
rect 16168 2688 16176 2752
rect 16240 2688 16256 2752
rect 16320 2688 16336 2752
rect 16400 2688 16416 2752
rect 16480 2688 16496 2752
rect 16560 2688 16568 2752
rect 14043 2548 14109 2549
rect 14043 2484 14044 2548
rect 14108 2484 14109 2548
rect 14043 2483 14109 2484
rect 10908 2144 10916 2208
rect 10980 2144 10996 2208
rect 11060 2144 11076 2208
rect 11140 2144 11156 2208
rect 11220 2144 11236 2208
rect 11300 2144 11308 2208
rect 10908 2128 11308 2144
rect 16168 2128 16568 2688
rect 16908 32672 17308 32688
rect 16908 32608 16916 32672
rect 16980 32608 16996 32672
rect 17060 32608 17076 32672
rect 17140 32608 17156 32672
rect 17220 32608 17236 32672
rect 17300 32608 17308 32672
rect 16908 31584 17308 32608
rect 16908 31520 16916 31584
rect 16980 31520 16996 31584
rect 17060 31520 17076 31584
rect 17140 31520 17156 31584
rect 17220 31520 17236 31584
rect 17300 31520 17308 31584
rect 16908 30496 17308 31520
rect 16908 30432 16916 30496
rect 16980 30432 16996 30496
rect 17060 30432 17076 30496
rect 17140 30432 17156 30496
rect 17220 30432 17236 30496
rect 17300 30432 17308 30496
rect 16908 30364 17308 30432
rect 16908 30128 16990 30364
rect 17226 30128 17308 30364
rect 16908 29408 17308 30128
rect 16908 29344 16916 29408
rect 16980 29344 16996 29408
rect 17060 29344 17076 29408
rect 17140 29344 17156 29408
rect 17220 29344 17236 29408
rect 17300 29344 17308 29408
rect 16908 28320 17308 29344
rect 16908 28256 16916 28320
rect 16980 28256 16996 28320
rect 17060 28256 17076 28320
rect 17140 28256 17156 28320
rect 17220 28256 17236 28320
rect 17300 28256 17308 28320
rect 16908 27232 17308 28256
rect 16908 27168 16916 27232
rect 16980 27168 16996 27232
rect 17060 27168 17076 27232
rect 17140 27168 17156 27232
rect 17220 27168 17236 27232
rect 17300 27168 17308 27232
rect 16908 26144 17308 27168
rect 16908 26080 16916 26144
rect 16980 26080 16996 26144
rect 17060 26080 17076 26144
rect 17140 26080 17156 26144
rect 17220 26080 17236 26144
rect 17300 26080 17308 26144
rect 16908 25056 17308 26080
rect 16908 24992 16916 25056
rect 16980 24992 16996 25056
rect 17060 24992 17076 25056
rect 17140 24992 17156 25056
rect 17220 24992 17236 25056
rect 17300 24992 17308 25056
rect 16908 24364 17308 24992
rect 16908 24128 16990 24364
rect 17226 24128 17308 24364
rect 16908 23968 17308 24128
rect 16908 23904 16916 23968
rect 16980 23904 16996 23968
rect 17060 23904 17076 23968
rect 17140 23904 17156 23968
rect 17220 23904 17236 23968
rect 17300 23904 17308 23968
rect 16908 22880 17308 23904
rect 16908 22816 16916 22880
rect 16980 22816 16996 22880
rect 17060 22816 17076 22880
rect 17140 22816 17156 22880
rect 17220 22816 17236 22880
rect 17300 22816 17308 22880
rect 16908 21792 17308 22816
rect 16908 21728 16916 21792
rect 16980 21728 16996 21792
rect 17060 21728 17076 21792
rect 17140 21728 17156 21792
rect 17220 21728 17236 21792
rect 17300 21728 17308 21792
rect 16908 20704 17308 21728
rect 22168 32128 22568 32688
rect 22168 32064 22176 32128
rect 22240 32064 22256 32128
rect 22320 32064 22336 32128
rect 22400 32064 22416 32128
rect 22480 32064 22496 32128
rect 22560 32064 22568 32128
rect 22168 31040 22568 32064
rect 22168 30976 22176 31040
rect 22240 30976 22256 31040
rect 22320 30976 22336 31040
rect 22400 30976 22416 31040
rect 22480 30976 22496 31040
rect 22560 30976 22568 31040
rect 22168 29952 22568 30976
rect 22168 29888 22176 29952
rect 22240 29888 22256 29952
rect 22320 29888 22336 29952
rect 22400 29888 22416 29952
rect 22480 29888 22496 29952
rect 22560 29888 22568 29952
rect 22168 29624 22568 29888
rect 22168 29388 22250 29624
rect 22486 29388 22568 29624
rect 22168 28864 22568 29388
rect 22168 28800 22176 28864
rect 22240 28800 22256 28864
rect 22320 28800 22336 28864
rect 22400 28800 22416 28864
rect 22480 28800 22496 28864
rect 22560 28800 22568 28864
rect 22168 27776 22568 28800
rect 22168 27712 22176 27776
rect 22240 27712 22256 27776
rect 22320 27712 22336 27776
rect 22400 27712 22416 27776
rect 22480 27712 22496 27776
rect 22560 27712 22568 27776
rect 22168 26688 22568 27712
rect 22168 26624 22176 26688
rect 22240 26624 22256 26688
rect 22320 26624 22336 26688
rect 22400 26624 22416 26688
rect 22480 26624 22496 26688
rect 22560 26624 22568 26688
rect 22168 25600 22568 26624
rect 22168 25536 22176 25600
rect 22240 25536 22256 25600
rect 22320 25536 22336 25600
rect 22400 25536 22416 25600
rect 22480 25536 22496 25600
rect 22560 25536 22568 25600
rect 22168 24512 22568 25536
rect 22168 24448 22176 24512
rect 22240 24448 22256 24512
rect 22320 24448 22336 24512
rect 22400 24448 22416 24512
rect 22480 24448 22496 24512
rect 22560 24448 22568 24512
rect 22168 23624 22568 24448
rect 22168 23424 22250 23624
rect 22486 23424 22568 23624
rect 22168 23360 22176 23424
rect 22240 23388 22250 23424
rect 22486 23388 22496 23424
rect 22240 23360 22256 23388
rect 22320 23360 22336 23388
rect 22400 23360 22416 23388
rect 22480 23360 22496 23388
rect 22560 23360 22568 23424
rect 22168 22336 22568 23360
rect 22168 22272 22176 22336
rect 22240 22272 22256 22336
rect 22320 22272 22336 22336
rect 22400 22272 22416 22336
rect 22480 22272 22496 22336
rect 22560 22272 22568 22336
rect 22168 21248 22568 22272
rect 22168 21184 22176 21248
rect 22240 21184 22256 21248
rect 22320 21184 22336 21248
rect 22400 21184 22416 21248
rect 22480 21184 22496 21248
rect 22560 21184 22568 21248
rect 20667 20772 20733 20773
rect 20667 20708 20668 20772
rect 20732 20708 20733 20772
rect 20667 20707 20733 20708
rect 16908 20640 16916 20704
rect 16980 20640 16996 20704
rect 17060 20640 17076 20704
rect 17140 20640 17156 20704
rect 17220 20640 17236 20704
rect 17300 20640 17308 20704
rect 16908 19616 17308 20640
rect 16908 19552 16916 19616
rect 16980 19552 16996 19616
rect 17060 19552 17076 19616
rect 17140 19552 17156 19616
rect 17220 19552 17236 19616
rect 17300 19552 17308 19616
rect 16908 18528 17308 19552
rect 16908 18464 16916 18528
rect 16980 18464 16996 18528
rect 17060 18464 17076 18528
rect 17140 18464 17156 18528
rect 17220 18464 17236 18528
rect 17300 18464 17308 18528
rect 16908 18364 17308 18464
rect 16908 18128 16990 18364
rect 17226 18128 17308 18364
rect 16908 17440 17308 18128
rect 20670 17509 20730 20707
rect 22168 20160 22568 21184
rect 22168 20096 22176 20160
rect 22240 20096 22256 20160
rect 22320 20096 22336 20160
rect 22400 20096 22416 20160
rect 22480 20096 22496 20160
rect 22560 20096 22568 20160
rect 22168 19072 22568 20096
rect 22168 19008 22176 19072
rect 22240 19008 22256 19072
rect 22320 19008 22336 19072
rect 22400 19008 22416 19072
rect 22480 19008 22496 19072
rect 22560 19008 22568 19072
rect 22168 17984 22568 19008
rect 22168 17920 22176 17984
rect 22240 17920 22256 17984
rect 22320 17920 22336 17984
rect 22400 17920 22416 17984
rect 22480 17920 22496 17984
rect 22560 17920 22568 17984
rect 22168 17624 22568 17920
rect 19379 17508 19445 17509
rect 19379 17444 19380 17508
rect 19444 17444 19445 17508
rect 19379 17443 19445 17444
rect 20667 17508 20733 17509
rect 20667 17444 20668 17508
rect 20732 17444 20733 17508
rect 20667 17443 20733 17444
rect 16908 17376 16916 17440
rect 16980 17376 16996 17440
rect 17060 17376 17076 17440
rect 17140 17376 17156 17440
rect 17220 17376 17236 17440
rect 17300 17376 17308 17440
rect 16908 16352 17308 17376
rect 16908 16288 16916 16352
rect 16980 16288 16996 16352
rect 17060 16288 17076 16352
rect 17140 16288 17156 16352
rect 17220 16288 17236 16352
rect 17300 16288 17308 16352
rect 16908 15264 17308 16288
rect 16908 15200 16916 15264
rect 16980 15200 16996 15264
rect 17060 15200 17076 15264
rect 17140 15200 17156 15264
rect 17220 15200 17236 15264
rect 17300 15200 17308 15264
rect 16908 14176 17308 15200
rect 16908 14112 16916 14176
rect 16980 14112 16996 14176
rect 17060 14112 17076 14176
rect 17140 14112 17156 14176
rect 17220 14112 17236 14176
rect 17300 14112 17308 14176
rect 16908 13088 17308 14112
rect 16908 13024 16916 13088
rect 16980 13024 16996 13088
rect 17060 13024 17076 13088
rect 17140 13024 17156 13088
rect 17220 13024 17236 13088
rect 17300 13024 17308 13088
rect 16908 12364 17308 13024
rect 19382 12749 19442 17443
rect 22168 17388 22250 17624
rect 22486 17388 22568 17624
rect 22168 16896 22568 17388
rect 22168 16832 22176 16896
rect 22240 16832 22256 16896
rect 22320 16832 22336 16896
rect 22400 16832 22416 16896
rect 22480 16832 22496 16896
rect 22560 16832 22568 16896
rect 22168 15808 22568 16832
rect 22168 15744 22176 15808
rect 22240 15744 22256 15808
rect 22320 15744 22336 15808
rect 22400 15744 22416 15808
rect 22480 15744 22496 15808
rect 22560 15744 22568 15808
rect 22168 14720 22568 15744
rect 22168 14656 22176 14720
rect 22240 14656 22256 14720
rect 22320 14656 22336 14720
rect 22400 14656 22416 14720
rect 22480 14656 22496 14720
rect 22560 14656 22568 14720
rect 22168 13632 22568 14656
rect 22168 13568 22176 13632
rect 22240 13568 22256 13632
rect 22320 13568 22336 13632
rect 22400 13568 22416 13632
rect 22480 13568 22496 13632
rect 22560 13568 22568 13632
rect 19379 12748 19445 12749
rect 19379 12684 19380 12748
rect 19444 12684 19445 12748
rect 19379 12683 19445 12684
rect 16908 12128 16990 12364
rect 17226 12128 17308 12364
rect 16908 12000 17308 12128
rect 16908 11936 16916 12000
rect 16980 11936 16996 12000
rect 17060 11936 17076 12000
rect 17140 11936 17156 12000
rect 17220 11936 17236 12000
rect 17300 11936 17308 12000
rect 16908 10912 17308 11936
rect 16908 10848 16916 10912
rect 16980 10848 16996 10912
rect 17060 10848 17076 10912
rect 17140 10848 17156 10912
rect 17220 10848 17236 10912
rect 17300 10848 17308 10912
rect 16908 9824 17308 10848
rect 16908 9760 16916 9824
rect 16980 9760 16996 9824
rect 17060 9760 17076 9824
rect 17140 9760 17156 9824
rect 17220 9760 17236 9824
rect 17300 9760 17308 9824
rect 16908 8736 17308 9760
rect 16908 8672 16916 8736
rect 16980 8672 16996 8736
rect 17060 8672 17076 8736
rect 17140 8672 17156 8736
rect 17220 8672 17236 8736
rect 17300 8672 17308 8736
rect 16908 7648 17308 8672
rect 16908 7584 16916 7648
rect 16980 7584 16996 7648
rect 17060 7584 17076 7648
rect 17140 7584 17156 7648
rect 17220 7584 17236 7648
rect 17300 7584 17308 7648
rect 16908 6560 17308 7584
rect 16908 6496 16916 6560
rect 16980 6496 16996 6560
rect 17060 6496 17076 6560
rect 17140 6496 17156 6560
rect 17220 6496 17236 6560
rect 17300 6496 17308 6560
rect 16908 6364 17308 6496
rect 16908 6128 16990 6364
rect 17226 6128 17308 6364
rect 16908 5472 17308 6128
rect 16908 5408 16916 5472
rect 16980 5408 16996 5472
rect 17060 5408 17076 5472
rect 17140 5408 17156 5472
rect 17220 5408 17236 5472
rect 17300 5408 17308 5472
rect 16908 4384 17308 5408
rect 16908 4320 16916 4384
rect 16980 4320 16996 4384
rect 17060 4320 17076 4384
rect 17140 4320 17156 4384
rect 17220 4320 17236 4384
rect 17300 4320 17308 4384
rect 16908 3296 17308 4320
rect 16908 3232 16916 3296
rect 16980 3232 16996 3296
rect 17060 3232 17076 3296
rect 17140 3232 17156 3296
rect 17220 3232 17236 3296
rect 17300 3232 17308 3296
rect 16908 2208 17308 3232
rect 16908 2144 16916 2208
rect 16980 2144 16996 2208
rect 17060 2144 17076 2208
rect 17140 2144 17156 2208
rect 17220 2144 17236 2208
rect 17300 2144 17308 2208
rect 16908 2128 17308 2144
rect 22168 12544 22568 13568
rect 22168 12480 22176 12544
rect 22240 12480 22256 12544
rect 22320 12480 22336 12544
rect 22400 12480 22416 12544
rect 22480 12480 22496 12544
rect 22560 12480 22568 12544
rect 22168 11624 22568 12480
rect 22168 11456 22250 11624
rect 22486 11456 22568 11624
rect 22168 11392 22176 11456
rect 22240 11392 22250 11456
rect 22486 11392 22496 11456
rect 22560 11392 22568 11456
rect 22168 11388 22250 11392
rect 22486 11388 22568 11392
rect 22168 10368 22568 11388
rect 22168 10304 22176 10368
rect 22240 10304 22256 10368
rect 22320 10304 22336 10368
rect 22400 10304 22416 10368
rect 22480 10304 22496 10368
rect 22560 10304 22568 10368
rect 22168 9280 22568 10304
rect 22168 9216 22176 9280
rect 22240 9216 22256 9280
rect 22320 9216 22336 9280
rect 22400 9216 22416 9280
rect 22480 9216 22496 9280
rect 22560 9216 22568 9280
rect 22168 8192 22568 9216
rect 22168 8128 22176 8192
rect 22240 8128 22256 8192
rect 22320 8128 22336 8192
rect 22400 8128 22416 8192
rect 22480 8128 22496 8192
rect 22560 8128 22568 8192
rect 22168 7104 22568 8128
rect 22168 7040 22176 7104
rect 22240 7040 22256 7104
rect 22320 7040 22336 7104
rect 22400 7040 22416 7104
rect 22480 7040 22496 7104
rect 22560 7040 22568 7104
rect 22168 6016 22568 7040
rect 22168 5952 22176 6016
rect 22240 5952 22256 6016
rect 22320 5952 22336 6016
rect 22400 5952 22416 6016
rect 22480 5952 22496 6016
rect 22560 5952 22568 6016
rect 22168 5624 22568 5952
rect 22168 5388 22250 5624
rect 22486 5388 22568 5624
rect 22168 4928 22568 5388
rect 22168 4864 22176 4928
rect 22240 4864 22256 4928
rect 22320 4864 22336 4928
rect 22400 4864 22416 4928
rect 22480 4864 22496 4928
rect 22560 4864 22568 4928
rect 22168 3840 22568 4864
rect 22168 3776 22176 3840
rect 22240 3776 22256 3840
rect 22320 3776 22336 3840
rect 22400 3776 22416 3840
rect 22480 3776 22496 3840
rect 22560 3776 22568 3840
rect 22168 2752 22568 3776
rect 22168 2688 22176 2752
rect 22240 2688 22256 2752
rect 22320 2688 22336 2752
rect 22400 2688 22416 2752
rect 22480 2688 22496 2752
rect 22560 2688 22568 2752
rect 22168 2128 22568 2688
rect 22908 32672 23308 32688
rect 22908 32608 22916 32672
rect 22980 32608 22996 32672
rect 23060 32608 23076 32672
rect 23140 32608 23156 32672
rect 23220 32608 23236 32672
rect 23300 32608 23308 32672
rect 22908 31584 23308 32608
rect 28168 32128 28568 32688
rect 28168 32064 28176 32128
rect 28240 32064 28256 32128
rect 28320 32064 28336 32128
rect 28400 32064 28416 32128
rect 28480 32064 28496 32128
rect 28560 32064 28568 32128
rect 27843 31924 27909 31925
rect 27843 31860 27844 31924
rect 27908 31860 27909 31924
rect 27843 31859 27909 31860
rect 22908 31520 22916 31584
rect 22980 31520 22996 31584
rect 23060 31520 23076 31584
rect 23140 31520 23156 31584
rect 23220 31520 23236 31584
rect 23300 31520 23308 31584
rect 22908 30496 23308 31520
rect 22908 30432 22916 30496
rect 22980 30432 22996 30496
rect 23060 30432 23076 30496
rect 23140 30432 23156 30496
rect 23220 30432 23236 30496
rect 23300 30432 23308 30496
rect 22908 30364 23308 30432
rect 22908 30128 22990 30364
rect 23226 30128 23308 30364
rect 22908 29408 23308 30128
rect 22908 29344 22916 29408
rect 22980 29344 22996 29408
rect 23060 29344 23076 29408
rect 23140 29344 23156 29408
rect 23220 29344 23236 29408
rect 23300 29344 23308 29408
rect 22908 28320 23308 29344
rect 22908 28256 22916 28320
rect 22980 28256 22996 28320
rect 23060 28256 23076 28320
rect 23140 28256 23156 28320
rect 23220 28256 23236 28320
rect 23300 28256 23308 28320
rect 22908 27232 23308 28256
rect 22908 27168 22916 27232
rect 22980 27168 22996 27232
rect 23060 27168 23076 27232
rect 23140 27168 23156 27232
rect 23220 27168 23236 27232
rect 23300 27168 23308 27232
rect 22908 26144 23308 27168
rect 22908 26080 22916 26144
rect 22980 26080 22996 26144
rect 23060 26080 23076 26144
rect 23140 26080 23156 26144
rect 23220 26080 23236 26144
rect 23300 26080 23308 26144
rect 22908 25056 23308 26080
rect 22908 24992 22916 25056
rect 22980 24992 22996 25056
rect 23060 24992 23076 25056
rect 23140 24992 23156 25056
rect 23220 24992 23236 25056
rect 23300 24992 23308 25056
rect 22908 24364 23308 24992
rect 22908 24128 22990 24364
rect 23226 24128 23308 24364
rect 22908 23968 23308 24128
rect 22908 23904 22916 23968
rect 22980 23904 22996 23968
rect 23060 23904 23076 23968
rect 23140 23904 23156 23968
rect 23220 23904 23236 23968
rect 23300 23904 23308 23968
rect 22908 22880 23308 23904
rect 22908 22816 22916 22880
rect 22980 22816 22996 22880
rect 23060 22816 23076 22880
rect 23140 22816 23156 22880
rect 23220 22816 23236 22880
rect 23300 22816 23308 22880
rect 22908 21792 23308 22816
rect 22908 21728 22916 21792
rect 22980 21728 22996 21792
rect 23060 21728 23076 21792
rect 23140 21728 23156 21792
rect 23220 21728 23236 21792
rect 23300 21728 23308 21792
rect 22908 20704 23308 21728
rect 22908 20640 22916 20704
rect 22980 20640 22996 20704
rect 23060 20640 23076 20704
rect 23140 20640 23156 20704
rect 23220 20640 23236 20704
rect 23300 20640 23308 20704
rect 22908 19616 23308 20640
rect 22908 19552 22916 19616
rect 22980 19552 22996 19616
rect 23060 19552 23076 19616
rect 23140 19552 23156 19616
rect 23220 19552 23236 19616
rect 23300 19552 23308 19616
rect 22908 18528 23308 19552
rect 22908 18464 22916 18528
rect 22980 18464 22996 18528
rect 23060 18464 23076 18528
rect 23140 18464 23156 18528
rect 23220 18464 23236 18528
rect 23300 18464 23308 18528
rect 22908 18364 23308 18464
rect 22908 18128 22990 18364
rect 23226 18128 23308 18364
rect 22908 17440 23308 18128
rect 27846 17645 27906 31859
rect 28168 31040 28568 32064
rect 28168 30976 28176 31040
rect 28240 30976 28256 31040
rect 28320 30976 28336 31040
rect 28400 30976 28416 31040
rect 28480 30976 28496 31040
rect 28560 30976 28568 31040
rect 28168 29952 28568 30976
rect 28168 29888 28176 29952
rect 28240 29888 28256 29952
rect 28320 29888 28336 29952
rect 28400 29888 28416 29952
rect 28480 29888 28496 29952
rect 28560 29888 28568 29952
rect 28168 29624 28568 29888
rect 28168 29388 28250 29624
rect 28486 29388 28568 29624
rect 28168 28864 28568 29388
rect 28168 28800 28176 28864
rect 28240 28800 28256 28864
rect 28320 28800 28336 28864
rect 28400 28800 28416 28864
rect 28480 28800 28496 28864
rect 28560 28800 28568 28864
rect 28168 27776 28568 28800
rect 28168 27712 28176 27776
rect 28240 27712 28256 27776
rect 28320 27712 28336 27776
rect 28400 27712 28416 27776
rect 28480 27712 28496 27776
rect 28560 27712 28568 27776
rect 28168 26688 28568 27712
rect 28168 26624 28176 26688
rect 28240 26624 28256 26688
rect 28320 26624 28336 26688
rect 28400 26624 28416 26688
rect 28480 26624 28496 26688
rect 28560 26624 28568 26688
rect 28168 25600 28568 26624
rect 28168 25536 28176 25600
rect 28240 25536 28256 25600
rect 28320 25536 28336 25600
rect 28400 25536 28416 25600
rect 28480 25536 28496 25600
rect 28560 25536 28568 25600
rect 28168 24512 28568 25536
rect 28168 24448 28176 24512
rect 28240 24448 28256 24512
rect 28320 24448 28336 24512
rect 28400 24448 28416 24512
rect 28480 24448 28496 24512
rect 28560 24448 28568 24512
rect 28168 23624 28568 24448
rect 28168 23424 28250 23624
rect 28486 23424 28568 23624
rect 28168 23360 28176 23424
rect 28240 23388 28250 23424
rect 28486 23388 28496 23424
rect 28240 23360 28256 23388
rect 28320 23360 28336 23388
rect 28400 23360 28416 23388
rect 28480 23360 28496 23388
rect 28560 23360 28568 23424
rect 28168 22336 28568 23360
rect 28168 22272 28176 22336
rect 28240 22272 28256 22336
rect 28320 22272 28336 22336
rect 28400 22272 28416 22336
rect 28480 22272 28496 22336
rect 28560 22272 28568 22336
rect 28168 21248 28568 22272
rect 28168 21184 28176 21248
rect 28240 21184 28256 21248
rect 28320 21184 28336 21248
rect 28400 21184 28416 21248
rect 28480 21184 28496 21248
rect 28560 21184 28568 21248
rect 28168 20160 28568 21184
rect 28168 20096 28176 20160
rect 28240 20096 28256 20160
rect 28320 20096 28336 20160
rect 28400 20096 28416 20160
rect 28480 20096 28496 20160
rect 28560 20096 28568 20160
rect 28168 19072 28568 20096
rect 28168 19008 28176 19072
rect 28240 19008 28256 19072
rect 28320 19008 28336 19072
rect 28400 19008 28416 19072
rect 28480 19008 28496 19072
rect 28560 19008 28568 19072
rect 28168 17984 28568 19008
rect 28168 17920 28176 17984
rect 28240 17920 28256 17984
rect 28320 17920 28336 17984
rect 28400 17920 28416 17984
rect 28480 17920 28496 17984
rect 28560 17920 28568 17984
rect 27843 17644 27909 17645
rect 27843 17580 27844 17644
rect 27908 17580 27909 17644
rect 27843 17579 27909 17580
rect 28168 17624 28568 17920
rect 22908 17376 22916 17440
rect 22980 17376 22996 17440
rect 23060 17376 23076 17440
rect 23140 17376 23156 17440
rect 23220 17376 23236 17440
rect 23300 17376 23308 17440
rect 22908 16352 23308 17376
rect 22908 16288 22916 16352
rect 22980 16288 22996 16352
rect 23060 16288 23076 16352
rect 23140 16288 23156 16352
rect 23220 16288 23236 16352
rect 23300 16288 23308 16352
rect 22908 15264 23308 16288
rect 22908 15200 22916 15264
rect 22980 15200 22996 15264
rect 23060 15200 23076 15264
rect 23140 15200 23156 15264
rect 23220 15200 23236 15264
rect 23300 15200 23308 15264
rect 22908 14176 23308 15200
rect 22908 14112 22916 14176
rect 22980 14112 22996 14176
rect 23060 14112 23076 14176
rect 23140 14112 23156 14176
rect 23220 14112 23236 14176
rect 23300 14112 23308 14176
rect 22908 13088 23308 14112
rect 22908 13024 22916 13088
rect 22980 13024 22996 13088
rect 23060 13024 23076 13088
rect 23140 13024 23156 13088
rect 23220 13024 23236 13088
rect 23300 13024 23308 13088
rect 22908 12364 23308 13024
rect 22908 12128 22990 12364
rect 23226 12128 23308 12364
rect 22908 12000 23308 12128
rect 22908 11936 22916 12000
rect 22980 11936 22996 12000
rect 23060 11936 23076 12000
rect 23140 11936 23156 12000
rect 23220 11936 23236 12000
rect 23300 11936 23308 12000
rect 22908 10912 23308 11936
rect 22908 10848 22916 10912
rect 22980 10848 22996 10912
rect 23060 10848 23076 10912
rect 23140 10848 23156 10912
rect 23220 10848 23236 10912
rect 23300 10848 23308 10912
rect 22908 9824 23308 10848
rect 22908 9760 22916 9824
rect 22980 9760 22996 9824
rect 23060 9760 23076 9824
rect 23140 9760 23156 9824
rect 23220 9760 23236 9824
rect 23300 9760 23308 9824
rect 22908 8736 23308 9760
rect 22908 8672 22916 8736
rect 22980 8672 22996 8736
rect 23060 8672 23076 8736
rect 23140 8672 23156 8736
rect 23220 8672 23236 8736
rect 23300 8672 23308 8736
rect 22908 7648 23308 8672
rect 22908 7584 22916 7648
rect 22980 7584 22996 7648
rect 23060 7584 23076 7648
rect 23140 7584 23156 7648
rect 23220 7584 23236 7648
rect 23300 7584 23308 7648
rect 22908 6560 23308 7584
rect 22908 6496 22916 6560
rect 22980 6496 22996 6560
rect 23060 6496 23076 6560
rect 23140 6496 23156 6560
rect 23220 6496 23236 6560
rect 23300 6496 23308 6560
rect 22908 6364 23308 6496
rect 22908 6128 22990 6364
rect 23226 6128 23308 6364
rect 22908 5472 23308 6128
rect 22908 5408 22916 5472
rect 22980 5408 22996 5472
rect 23060 5408 23076 5472
rect 23140 5408 23156 5472
rect 23220 5408 23236 5472
rect 23300 5408 23308 5472
rect 22908 4384 23308 5408
rect 22908 4320 22916 4384
rect 22980 4320 22996 4384
rect 23060 4320 23076 4384
rect 23140 4320 23156 4384
rect 23220 4320 23236 4384
rect 23300 4320 23308 4384
rect 22908 3296 23308 4320
rect 22908 3232 22916 3296
rect 22980 3232 22996 3296
rect 23060 3232 23076 3296
rect 23140 3232 23156 3296
rect 23220 3232 23236 3296
rect 23300 3232 23308 3296
rect 22908 2208 23308 3232
rect 22908 2144 22916 2208
rect 22980 2144 22996 2208
rect 23060 2144 23076 2208
rect 23140 2144 23156 2208
rect 23220 2144 23236 2208
rect 23300 2144 23308 2208
rect 22908 2128 23308 2144
rect 28168 17388 28250 17624
rect 28486 17388 28568 17624
rect 28168 16896 28568 17388
rect 28168 16832 28176 16896
rect 28240 16832 28256 16896
rect 28320 16832 28336 16896
rect 28400 16832 28416 16896
rect 28480 16832 28496 16896
rect 28560 16832 28568 16896
rect 28168 15808 28568 16832
rect 28168 15744 28176 15808
rect 28240 15744 28256 15808
rect 28320 15744 28336 15808
rect 28400 15744 28416 15808
rect 28480 15744 28496 15808
rect 28560 15744 28568 15808
rect 28168 14720 28568 15744
rect 28168 14656 28176 14720
rect 28240 14656 28256 14720
rect 28320 14656 28336 14720
rect 28400 14656 28416 14720
rect 28480 14656 28496 14720
rect 28560 14656 28568 14720
rect 28168 13632 28568 14656
rect 28168 13568 28176 13632
rect 28240 13568 28256 13632
rect 28320 13568 28336 13632
rect 28400 13568 28416 13632
rect 28480 13568 28496 13632
rect 28560 13568 28568 13632
rect 28168 12544 28568 13568
rect 28168 12480 28176 12544
rect 28240 12480 28256 12544
rect 28320 12480 28336 12544
rect 28400 12480 28416 12544
rect 28480 12480 28496 12544
rect 28560 12480 28568 12544
rect 28168 11624 28568 12480
rect 28168 11456 28250 11624
rect 28486 11456 28568 11624
rect 28168 11392 28176 11456
rect 28240 11392 28250 11456
rect 28486 11392 28496 11456
rect 28560 11392 28568 11456
rect 28168 11388 28250 11392
rect 28486 11388 28568 11392
rect 28168 10368 28568 11388
rect 28168 10304 28176 10368
rect 28240 10304 28256 10368
rect 28320 10304 28336 10368
rect 28400 10304 28416 10368
rect 28480 10304 28496 10368
rect 28560 10304 28568 10368
rect 28168 9280 28568 10304
rect 28168 9216 28176 9280
rect 28240 9216 28256 9280
rect 28320 9216 28336 9280
rect 28400 9216 28416 9280
rect 28480 9216 28496 9280
rect 28560 9216 28568 9280
rect 28168 8192 28568 9216
rect 28168 8128 28176 8192
rect 28240 8128 28256 8192
rect 28320 8128 28336 8192
rect 28400 8128 28416 8192
rect 28480 8128 28496 8192
rect 28560 8128 28568 8192
rect 28168 7104 28568 8128
rect 28168 7040 28176 7104
rect 28240 7040 28256 7104
rect 28320 7040 28336 7104
rect 28400 7040 28416 7104
rect 28480 7040 28496 7104
rect 28560 7040 28568 7104
rect 28168 6016 28568 7040
rect 28168 5952 28176 6016
rect 28240 5952 28256 6016
rect 28320 5952 28336 6016
rect 28400 5952 28416 6016
rect 28480 5952 28496 6016
rect 28560 5952 28568 6016
rect 28168 5624 28568 5952
rect 28168 5388 28250 5624
rect 28486 5388 28568 5624
rect 28168 4928 28568 5388
rect 28168 4864 28176 4928
rect 28240 4864 28256 4928
rect 28320 4864 28336 4928
rect 28400 4864 28416 4928
rect 28480 4864 28496 4928
rect 28560 4864 28568 4928
rect 28168 3840 28568 4864
rect 28168 3776 28176 3840
rect 28240 3776 28256 3840
rect 28320 3776 28336 3840
rect 28400 3776 28416 3840
rect 28480 3776 28496 3840
rect 28560 3776 28568 3840
rect 28168 2752 28568 3776
rect 28168 2688 28176 2752
rect 28240 2688 28256 2752
rect 28320 2688 28336 2752
rect 28400 2688 28416 2752
rect 28480 2688 28496 2752
rect 28560 2688 28568 2752
rect 28168 2128 28568 2688
rect 28908 32672 29308 32688
rect 28908 32608 28916 32672
rect 28980 32608 28996 32672
rect 29060 32608 29076 32672
rect 29140 32608 29156 32672
rect 29220 32608 29236 32672
rect 29300 32608 29308 32672
rect 28908 31584 29308 32608
rect 28908 31520 28916 31584
rect 28980 31520 28996 31584
rect 29060 31520 29076 31584
rect 29140 31520 29156 31584
rect 29220 31520 29236 31584
rect 29300 31520 29308 31584
rect 28908 30496 29308 31520
rect 28908 30432 28916 30496
rect 28980 30432 28996 30496
rect 29060 30432 29076 30496
rect 29140 30432 29156 30496
rect 29220 30432 29236 30496
rect 29300 30432 29308 30496
rect 28908 30364 29308 30432
rect 28908 30128 28990 30364
rect 29226 30128 29308 30364
rect 28908 29408 29308 30128
rect 28908 29344 28916 29408
rect 28980 29344 28996 29408
rect 29060 29344 29076 29408
rect 29140 29344 29156 29408
rect 29220 29344 29236 29408
rect 29300 29344 29308 29408
rect 28908 28320 29308 29344
rect 28908 28256 28916 28320
rect 28980 28256 28996 28320
rect 29060 28256 29076 28320
rect 29140 28256 29156 28320
rect 29220 28256 29236 28320
rect 29300 28256 29308 28320
rect 28908 27232 29308 28256
rect 28908 27168 28916 27232
rect 28980 27168 28996 27232
rect 29060 27168 29076 27232
rect 29140 27168 29156 27232
rect 29220 27168 29236 27232
rect 29300 27168 29308 27232
rect 28908 26144 29308 27168
rect 28908 26080 28916 26144
rect 28980 26080 28996 26144
rect 29060 26080 29076 26144
rect 29140 26080 29156 26144
rect 29220 26080 29236 26144
rect 29300 26080 29308 26144
rect 28908 25056 29308 26080
rect 28908 24992 28916 25056
rect 28980 24992 28996 25056
rect 29060 24992 29076 25056
rect 29140 24992 29156 25056
rect 29220 24992 29236 25056
rect 29300 24992 29308 25056
rect 28908 24364 29308 24992
rect 28908 24128 28990 24364
rect 29226 24128 29308 24364
rect 28908 23968 29308 24128
rect 28908 23904 28916 23968
rect 28980 23904 28996 23968
rect 29060 23904 29076 23968
rect 29140 23904 29156 23968
rect 29220 23904 29236 23968
rect 29300 23904 29308 23968
rect 28908 22880 29308 23904
rect 28908 22816 28916 22880
rect 28980 22816 28996 22880
rect 29060 22816 29076 22880
rect 29140 22816 29156 22880
rect 29220 22816 29236 22880
rect 29300 22816 29308 22880
rect 28908 21792 29308 22816
rect 28908 21728 28916 21792
rect 28980 21728 28996 21792
rect 29060 21728 29076 21792
rect 29140 21728 29156 21792
rect 29220 21728 29236 21792
rect 29300 21728 29308 21792
rect 28908 20704 29308 21728
rect 28908 20640 28916 20704
rect 28980 20640 28996 20704
rect 29060 20640 29076 20704
rect 29140 20640 29156 20704
rect 29220 20640 29236 20704
rect 29300 20640 29308 20704
rect 28908 19616 29308 20640
rect 28908 19552 28916 19616
rect 28980 19552 28996 19616
rect 29060 19552 29076 19616
rect 29140 19552 29156 19616
rect 29220 19552 29236 19616
rect 29300 19552 29308 19616
rect 28908 18528 29308 19552
rect 28908 18464 28916 18528
rect 28980 18464 28996 18528
rect 29060 18464 29076 18528
rect 29140 18464 29156 18528
rect 29220 18464 29236 18528
rect 29300 18464 29308 18528
rect 28908 18364 29308 18464
rect 28908 18128 28990 18364
rect 29226 18128 29308 18364
rect 28908 17440 29308 18128
rect 28908 17376 28916 17440
rect 28980 17376 28996 17440
rect 29060 17376 29076 17440
rect 29140 17376 29156 17440
rect 29220 17376 29236 17440
rect 29300 17376 29308 17440
rect 28908 16352 29308 17376
rect 28908 16288 28916 16352
rect 28980 16288 28996 16352
rect 29060 16288 29076 16352
rect 29140 16288 29156 16352
rect 29220 16288 29236 16352
rect 29300 16288 29308 16352
rect 28908 15264 29308 16288
rect 28908 15200 28916 15264
rect 28980 15200 28996 15264
rect 29060 15200 29076 15264
rect 29140 15200 29156 15264
rect 29220 15200 29236 15264
rect 29300 15200 29308 15264
rect 28908 14176 29308 15200
rect 28908 14112 28916 14176
rect 28980 14112 28996 14176
rect 29060 14112 29076 14176
rect 29140 14112 29156 14176
rect 29220 14112 29236 14176
rect 29300 14112 29308 14176
rect 28908 13088 29308 14112
rect 28908 13024 28916 13088
rect 28980 13024 28996 13088
rect 29060 13024 29076 13088
rect 29140 13024 29156 13088
rect 29220 13024 29236 13088
rect 29300 13024 29308 13088
rect 28908 12364 29308 13024
rect 28908 12128 28990 12364
rect 29226 12128 29308 12364
rect 28908 12000 29308 12128
rect 28908 11936 28916 12000
rect 28980 11936 28996 12000
rect 29060 11936 29076 12000
rect 29140 11936 29156 12000
rect 29220 11936 29236 12000
rect 29300 11936 29308 12000
rect 28908 10912 29308 11936
rect 28908 10848 28916 10912
rect 28980 10848 28996 10912
rect 29060 10848 29076 10912
rect 29140 10848 29156 10912
rect 29220 10848 29236 10912
rect 29300 10848 29308 10912
rect 28908 9824 29308 10848
rect 28908 9760 28916 9824
rect 28980 9760 28996 9824
rect 29060 9760 29076 9824
rect 29140 9760 29156 9824
rect 29220 9760 29236 9824
rect 29300 9760 29308 9824
rect 28908 8736 29308 9760
rect 28908 8672 28916 8736
rect 28980 8672 28996 8736
rect 29060 8672 29076 8736
rect 29140 8672 29156 8736
rect 29220 8672 29236 8736
rect 29300 8672 29308 8736
rect 28908 7648 29308 8672
rect 28908 7584 28916 7648
rect 28980 7584 28996 7648
rect 29060 7584 29076 7648
rect 29140 7584 29156 7648
rect 29220 7584 29236 7648
rect 29300 7584 29308 7648
rect 28908 6560 29308 7584
rect 28908 6496 28916 6560
rect 28980 6496 28996 6560
rect 29060 6496 29076 6560
rect 29140 6496 29156 6560
rect 29220 6496 29236 6560
rect 29300 6496 29308 6560
rect 28908 6364 29308 6496
rect 28908 6128 28990 6364
rect 29226 6128 29308 6364
rect 28908 5472 29308 6128
rect 28908 5408 28916 5472
rect 28980 5408 28996 5472
rect 29060 5408 29076 5472
rect 29140 5408 29156 5472
rect 29220 5408 29236 5472
rect 29300 5408 29308 5472
rect 28908 4384 29308 5408
rect 28908 4320 28916 4384
rect 28980 4320 28996 4384
rect 29060 4320 29076 4384
rect 29140 4320 29156 4384
rect 29220 4320 29236 4384
rect 29300 4320 29308 4384
rect 28908 3296 29308 4320
rect 28908 3232 28916 3296
rect 28980 3232 28996 3296
rect 29060 3232 29076 3296
rect 29140 3232 29156 3296
rect 29220 3232 29236 3296
rect 29300 3232 29308 3296
rect 28908 2208 29308 3232
rect 28908 2144 28916 2208
rect 28980 2144 28996 2208
rect 29060 2144 29076 2208
rect 29140 2144 29156 2208
rect 29220 2144 29236 2208
rect 29300 2144 29308 2208
rect 28908 2128 29308 2144
<< via4 >>
rect 4250 29388 4486 29624
rect 4250 23424 4486 23624
rect 4250 23388 4256 23424
rect 4256 23388 4320 23424
rect 4320 23388 4336 23424
rect 4336 23388 4400 23424
rect 4400 23388 4416 23424
rect 4416 23388 4480 23424
rect 4480 23388 4486 23424
rect 4250 17388 4486 17624
rect 4250 11456 4486 11624
rect 4250 11392 4256 11456
rect 4256 11392 4320 11456
rect 4320 11392 4336 11456
rect 4336 11392 4400 11456
rect 4400 11392 4416 11456
rect 4416 11392 4480 11456
rect 4480 11392 4486 11456
rect 4250 11388 4486 11392
rect 4250 5388 4486 5624
rect 4990 30128 5226 30364
rect 4990 24128 5226 24364
rect 4990 18128 5226 18364
rect 4990 12128 5226 12364
rect 10250 29388 10486 29624
rect 10250 23424 10486 23624
rect 10250 23388 10256 23424
rect 10256 23388 10320 23424
rect 10320 23388 10336 23424
rect 10336 23388 10400 23424
rect 10400 23388 10416 23424
rect 10416 23388 10480 23424
rect 10480 23388 10486 23424
rect 10250 17388 10486 17624
rect 10250 11456 10486 11624
rect 10250 11392 10256 11456
rect 10256 11392 10320 11456
rect 10320 11392 10336 11456
rect 10336 11392 10400 11456
rect 10400 11392 10416 11456
rect 10416 11392 10480 11456
rect 10480 11392 10486 11456
rect 10250 11388 10486 11392
rect 4990 6128 5226 6364
rect 10990 30128 11226 30364
rect 16250 29388 16486 29624
rect 10990 24128 11226 24364
rect 10990 18128 11226 18364
rect 10990 12128 11226 12364
rect 10250 5388 10486 5624
rect 10990 6128 11226 6364
rect 16250 23424 16486 23624
rect 16250 23388 16256 23424
rect 16256 23388 16320 23424
rect 16320 23388 16336 23424
rect 16336 23388 16400 23424
rect 16400 23388 16416 23424
rect 16416 23388 16480 23424
rect 16480 23388 16486 23424
rect 16250 17388 16486 17624
rect 16250 11456 16486 11624
rect 16250 11392 16256 11456
rect 16256 11392 16320 11456
rect 16320 11392 16336 11456
rect 16336 11392 16400 11456
rect 16400 11392 16416 11456
rect 16416 11392 16480 11456
rect 16480 11392 16486 11456
rect 16250 11388 16486 11392
rect 16250 5388 16486 5624
rect 16990 30128 17226 30364
rect 16990 24128 17226 24364
rect 22250 29388 22486 29624
rect 22250 23424 22486 23624
rect 22250 23388 22256 23424
rect 22256 23388 22320 23424
rect 22320 23388 22336 23424
rect 22336 23388 22400 23424
rect 22400 23388 22416 23424
rect 22416 23388 22480 23424
rect 22480 23388 22486 23424
rect 16990 18128 17226 18364
rect 22250 17388 22486 17624
rect 16990 12128 17226 12364
rect 16990 6128 17226 6364
rect 22250 11456 22486 11624
rect 22250 11392 22256 11456
rect 22256 11392 22320 11456
rect 22320 11392 22336 11456
rect 22336 11392 22400 11456
rect 22400 11392 22416 11456
rect 22416 11392 22480 11456
rect 22480 11392 22486 11456
rect 22250 11388 22486 11392
rect 22250 5388 22486 5624
rect 22990 30128 23226 30364
rect 22990 24128 23226 24364
rect 22990 18128 23226 18364
rect 28250 29388 28486 29624
rect 28250 23424 28486 23624
rect 28250 23388 28256 23424
rect 28256 23388 28320 23424
rect 28320 23388 28336 23424
rect 28336 23388 28400 23424
rect 28400 23388 28416 23424
rect 28416 23388 28480 23424
rect 28480 23388 28486 23424
rect 22990 12128 23226 12364
rect 22990 6128 23226 6364
rect 28250 17388 28486 17624
rect 28250 11456 28486 11624
rect 28250 11392 28256 11456
rect 28256 11392 28320 11456
rect 28320 11392 28336 11456
rect 28336 11392 28400 11456
rect 28400 11392 28416 11456
rect 28416 11392 28480 11456
rect 28480 11392 28486 11456
rect 28250 11388 28486 11392
rect 28250 5388 28486 5624
rect 28990 30128 29226 30364
rect 28990 24128 29226 24364
rect 28990 18128 29226 18364
rect 28990 12128 29226 12364
rect 28990 6128 29226 6364
<< metal5 >>
rect 1056 30364 31880 30446
rect 1056 30128 4990 30364
rect 5226 30128 10990 30364
rect 11226 30128 16990 30364
rect 17226 30128 22990 30364
rect 23226 30128 28990 30364
rect 29226 30128 31880 30364
rect 1056 30046 31880 30128
rect 1056 29624 31880 29706
rect 1056 29388 4250 29624
rect 4486 29388 10250 29624
rect 10486 29388 16250 29624
rect 16486 29388 22250 29624
rect 22486 29388 28250 29624
rect 28486 29388 31880 29624
rect 1056 29306 31880 29388
rect 1056 24364 31880 24446
rect 1056 24128 4990 24364
rect 5226 24128 10990 24364
rect 11226 24128 16990 24364
rect 17226 24128 22990 24364
rect 23226 24128 28990 24364
rect 29226 24128 31880 24364
rect 1056 24046 31880 24128
rect 1056 23624 31880 23706
rect 1056 23388 4250 23624
rect 4486 23388 10250 23624
rect 10486 23388 16250 23624
rect 16486 23388 22250 23624
rect 22486 23388 28250 23624
rect 28486 23388 31880 23624
rect 1056 23306 31880 23388
rect 1056 18364 31880 18446
rect 1056 18128 4990 18364
rect 5226 18128 10990 18364
rect 11226 18128 16990 18364
rect 17226 18128 22990 18364
rect 23226 18128 28990 18364
rect 29226 18128 31880 18364
rect 1056 18046 31880 18128
rect 1056 17624 31880 17706
rect 1056 17388 4250 17624
rect 4486 17388 10250 17624
rect 10486 17388 16250 17624
rect 16486 17388 22250 17624
rect 22486 17388 28250 17624
rect 28486 17388 31880 17624
rect 1056 17306 31880 17388
rect 1056 12364 31880 12446
rect 1056 12128 4990 12364
rect 5226 12128 10990 12364
rect 11226 12128 16990 12364
rect 17226 12128 22990 12364
rect 23226 12128 28990 12364
rect 29226 12128 31880 12364
rect 1056 12046 31880 12128
rect 1056 11624 31880 11706
rect 1056 11388 4250 11624
rect 4486 11388 10250 11624
rect 10486 11388 16250 11624
rect 16486 11388 22250 11624
rect 22486 11388 28250 11624
rect 28486 11388 31880 11624
rect 1056 11306 31880 11388
rect 1056 6364 31880 6446
rect 1056 6128 4990 6364
rect 5226 6128 10990 6364
rect 11226 6128 16990 6364
rect 17226 6128 22990 6364
rect 23226 6128 28990 6364
rect 29226 6128 31880 6364
rect 1056 6046 31880 6128
rect 1056 5624 31880 5706
rect 1056 5388 4250 5624
rect 4486 5388 10250 5624
rect 10486 5388 16250 5624
rect 16486 5388 22250 5624
rect 22486 5388 28250 5624
rect 28486 5388 31880 5624
rect 1056 5306 31880 5388
use sky130_fd_sc_hd__xnor2_1  _0489_
timestamp 0
transform 1 0 19228 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0490_
timestamp 0
transform 1 0 19872 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0491_
timestamp 0
transform 1 0 20148 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0492_
timestamp 0
transform 1 0 20332 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and4_2  _0493_
timestamp 0
transform 1 0 20700 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_4  _0494_
timestamp 0
transform 1 0 11592 0 -1 30464
box -38 -48 2062 592
use sky130_fd_sc_hd__a21boi_4  _0495_
timestamp 0
transform 1 0 12512 0 -1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__buf_2  _0496_
timestamp 0
transform 1 0 20424 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__and4b_1  _0497_
timestamp 0
transform 1 0 19412 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _0498_
timestamp 0
transform 1 0 19964 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0499_
timestamp 0
transform -1 0 19504 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0500_
timestamp 0
transform 1 0 14996 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _0501_
timestamp 0
transform 1 0 13892 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0502_
timestamp 0
transform 1 0 19780 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0503_
timestamp 0
transform 1 0 20240 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0504_
timestamp 0
transform -1 0 14444 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0505_
timestamp 0
transform 1 0 15088 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0506_
timestamp 0
transform 1 0 18768 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0507_
timestamp 0
transform 1 0 15272 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0508_
timestamp 0
transform 1 0 15548 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0509_
timestamp 0
transform 1 0 16192 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0510_
timestamp 0
transform -1 0 14720 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0511_
timestamp 0
transform -1 0 15180 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0512_
timestamp 0
transform -1 0 16376 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0513_
timestamp 0
transform -1 0 15824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0514_
timestamp 0
transform -1 0 16376 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0515_
timestamp 0
transform -1 0 14352 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _0516_
timestamp 0
transform 1 0 12972 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0517_
timestamp 0
transform 1 0 14536 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__and2_2  _0518_
timestamp 0
transform -1 0 17940 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0519_
timestamp 0
transform -1 0 16652 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0520_
timestamp 0
transform -1 0 15180 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0521_
timestamp 0
transform -1 0 17112 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _0522_
timestamp 0
transform 1 0 15640 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0523_
timestamp 0
transform -1 0 17388 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0524_
timestamp 0
transform -1 0 18400 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0525_
timestamp 0
transform 1 0 15456 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0526_
timestamp 0
transform -1 0 17756 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0527_
timestamp 0
transform -1 0 18124 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _0528_
timestamp 0
transform 1 0 17664 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0529_
timestamp 0
transform -1 0 12236 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__nor4b_1  _0530_
timestamp 0
transform -1 0 22908 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_4  _0531_
timestamp 0
transform -1 0 23000 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__nor4_1  _0532_
timestamp 0
transform 1 0 21252 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0533_
timestamp 0
transform -1 0 29256 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nor4b_1  _0534_
timestamp 0
transform -1 0 21896 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nor4b_1  _0535_
timestamp 0
transform -1 0 20792 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0536_
timestamp 0
transform 1 0 26036 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_4  _0537_
timestamp 0
transform 1 0 19504 0 -1 23936
box -38 -48 1050 592
use sky130_fd_sc_hd__and4bb_4  _0538_
timestamp 0
transform -1 0 20608 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__a22o_1  _0539_
timestamp 0
transform 1 0 26220 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_4  _0540_
timestamp 0
transform 1 0 20516 0 -1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__and4bb_4  _0541_
timestamp 0
transform -1 0 21804 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__a22o_1  _0542_
timestamp 0
transform 1 0 23920 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0543_
timestamp 0
transform 1 0 26956 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and4bb_4  _0544_
timestamp 0
transform 1 0 13892 0 -1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__and4b_4  _0545_
timestamp 0
transform 1 0 12788 0 -1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__and4b_4  _0546_
timestamp 0
transform 1 0 12788 0 1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__a22o_1  _0547_
timestamp 0
transform 1 0 5980 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0548_
timestamp 0
transform 1 0 7544 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _0549_
timestamp 0
transform -1 0 14076 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _0550_
timestamp 0
transform 1 0 13248 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _0551_
timestamp 0
transform 1 0 14076 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__and4bb_4  _0552_
timestamp 0
transform -1 0 13892 0 -1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__a22o_1  _0553_
timestamp 0
transform -1 0 9936 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0554_
timestamp 0
transform 1 0 8924 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or4_4  _0555_
timestamp 0
transform 1 0 14076 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0556_
timestamp 0
transform -1 0 11132 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _0557_
timestamp 0
transform -1 0 10396 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0558_
timestamp 0
transform 1 0 9660 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0559_
timestamp 0
transform 1 0 9292 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _0560_
timestamp 0
transform -1 0 29164 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0561_
timestamp 0
transform 1 0 25392 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0562_
timestamp 0
transform -1 0 27600 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0563_
timestamp 0
transform 1 0 24196 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0564_
timestamp 0
transform 1 0 25760 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0565_
timestamp 0
transform 1 0 5520 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0566_
timestamp 0
transform -1 0 8556 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0567_
timestamp 0
transform -1 0 10304 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0568_
timestamp 0
transform 1 0 9660 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0569_
timestamp 0
transform -1 0 12236 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _0570_
timestamp 0
transform -1 0 11776 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0571_
timestamp 0
transform -1 0 13248 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0572_
timestamp 0
transform 1 0 13248 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _0573_
timestamp 0
transform -1 0 29440 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0574_
timestamp 0
transform -1 0 26864 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0575_
timestamp 0
transform -1 0 26680 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0576_
timestamp 0
transform 1 0 23276 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0577_
timestamp 0
transform -1 0 26036 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0578_
timestamp 0
transform 1 0 5796 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0579_
timestamp 0
transform -1 0 9292 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0580_
timestamp 0
transform 1 0 7728 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0581_
timestamp 0
transform 1 0 8924 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0582_
timestamp 0
transform -1 0 11960 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _0583_
timestamp 0
transform -1 0 10488 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0584_
timestamp 0
transform 1 0 10488 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0585_
timestamp 0
transform -1 0 10304 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _0586_
timestamp 0
transform -1 0 27692 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0587_
timestamp 0
transform -1 0 23368 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0588_
timestamp 0
transform 1 0 19228 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0589_
timestamp 0
transform 1 0 20424 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0590_
timestamp 0
transform 1 0 21160 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0591_
timestamp 0
transform 1 0 5336 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0592_
timestamp 0
transform -1 0 15364 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0593_
timestamp 0
transform 1 0 12144 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0594_
timestamp 0
transform 1 0 13248 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0595_
timestamp 0
transform 1 0 15916 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _0596_
timestamp 0
transform 1 0 16008 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0597_
timestamp 0
transform -1 0 15456 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0598_
timestamp 0
transform -1 0 15364 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _0599_
timestamp 0
transform -1 0 21620 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0600_
timestamp 0
transform -1 0 21436 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0601_
timestamp 0
transform 1 0 18492 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0602_
timestamp 0
transform 1 0 18952 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0603_
timestamp 0
transform 1 0 19596 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0604_
timestamp 0
transform 1 0 4876 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0605_
timestamp 0
transform -1 0 8924 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0606_
timestamp 0
transform 1 0 8556 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0607_
timestamp 0
transform 1 0 9200 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0608_
timestamp 0
transform -1 0 11224 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _0609_
timestamp 0
transform 1 0 9936 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0610_
timestamp 0
transform 1 0 9384 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0611_
timestamp 0
transform 1 0 9108 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _0612_
timestamp 0
transform -1 0 24288 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0613_
timestamp 0
transform -1 0 23368 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0614_
timestamp 0
transform 1 0 21896 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0615_
timestamp 0
transform 1 0 21804 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0616_
timestamp 0
transform 1 0 22540 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0617_
timestamp 0
transform 1 0 5520 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0618_
timestamp 0
transform 1 0 7820 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0619_
timestamp 0
transform 1 0 8096 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0620_
timestamp 0
transform 1 0 9016 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0621_
timestamp 0
transform -1 0 11960 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _0622_
timestamp 0
transform 1 0 10856 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0623_
timestamp 0
transform 1 0 9660 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0624_
timestamp 0
transform 1 0 9476 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _0625_
timestamp 0
transform 1 0 30360 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0626_
timestamp 0
transform -1 0 26772 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0627_
timestamp 0
transform -1 0 26864 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0628_
timestamp 0
transform 1 0 25944 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0629_
timestamp 0
transform 1 0 26404 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0630_
timestamp 0
transform 1 0 7820 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0631_
timestamp 0
transform -1 0 14628 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0632_
timestamp 0
transform 1 0 13156 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0633_
timestamp 0
transform 1 0 13892 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0634_
timestamp 0
transform 1 0 16100 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _0635_
timestamp 0
transform 1 0 14628 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0636_
timestamp 0
transform 1 0 14076 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0637_
timestamp 0
transform 1 0 13064 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _0638_
timestamp 0
transform -1 0 30268 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0639_
timestamp 0
transform -1 0 25392 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0640_
timestamp 0
transform 1 0 19780 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0641_
timestamp 0
transform 1 0 20424 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0642_
timestamp 0
transform 1 0 21804 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0643_
timestamp 0
transform 1 0 4692 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0644_
timestamp 0
transform -1 0 16836 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0645_
timestamp 0
transform 1 0 12788 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0646_
timestamp 0
transform 1 0 13616 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0647_
timestamp 0
transform 1 0 15732 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _0648_
timestamp 0
transform 1 0 15640 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0649_
timestamp 0
transform 1 0 15456 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0650_
timestamp 0
transform -1 0 15640 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0651_
timestamp 0
transform -1 0 11132 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0652_
timestamp 0
transform 1 0 13524 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0653_
timestamp 0
transform 1 0 13800 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0654_
timestamp 0
transform -1 0 14536 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _0655_
timestamp 0
transform -1 0 13800 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0656_
timestamp 0
transform 1 0 13156 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0657_
timestamp 0
transform -1 0 19044 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0658_
timestamp 0
transform 1 0 19228 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  _0659_
timestamp 0
transform -1 0 17664 0 -1 30464
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_2  _0660_
timestamp 0
transform 1 0 16652 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0661_
timestamp 0
transform -1 0 13892 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0662_
timestamp 0
transform -1 0 10028 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0663_
timestamp 0
transform -1 0 10764 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0664_
timestamp 0
transform 1 0 16192 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0665_
timestamp 0
transform -1 0 11776 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0666_
timestamp 0
transform -1 0 14352 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0667_
timestamp 0
transform -1 0 11040 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0668_
timestamp 0
transform -1 0 13340 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0669_
timestamp 0
transform 1 0 14720 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0670_
timestamp 0
transform 1 0 19596 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0671_
timestamp 0
transform 1 0 19320 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0672_
timestamp 0
transform 1 0 18492 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0673_
timestamp 0
transform -1 0 17020 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0674_
timestamp 0
transform -1 0 18676 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0675_
timestamp 0
transform -1 0 19044 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0676_
timestamp 0
transform -1 0 19504 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0677_
timestamp 0
transform -1 0 17664 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0678_
timestamp 0
transform 1 0 16652 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0679_
timestamp 0
transform 1 0 14720 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _0680_
timestamp 0
transform -1 0 19044 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0681_
timestamp 0
transform 1 0 16652 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _0682_
timestamp 0
transform 1 0 14536 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _0683_
timestamp 0
transform -1 0 15272 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0684_
timestamp 0
transform 1 0 14904 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0685_
timestamp 0
transform -1 0 14628 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0686_
timestamp 0
transform 1 0 28612 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0687_
timestamp 0
transform -1 0 15180 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0688_
timestamp 0
transform 1 0 14628 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0689_
timestamp 0
transform 1 0 16560 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0690_
timestamp 0
transform 1 0 11868 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0691_
timestamp 0
transform -1 0 11408 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0692_
timestamp 0
transform 1 0 17112 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0693_
timestamp 0
transform 1 0 11500 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0694_
timestamp 0
transform 1 0 10672 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0695_
timestamp 0
transform 1 0 16928 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0696_
timestamp 0
transform 1 0 14444 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0697_
timestamp 0
transform -1 0 13340 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0698_
timestamp 0
transform 1 0 15088 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0699_
timestamp 0
transform 1 0 10488 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0700_
timestamp 0
transform 1 0 10212 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0701_
timestamp 0
transform 1 0 29072 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0702_
timestamp 0
transform 1 0 11500 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0703_
timestamp 0
transform 1 0 11132 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0704_
timestamp 0
transform 1 0 28060 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0705_
timestamp 0
transform 1 0 10580 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0706_
timestamp 0
transform 1 0 10396 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0707_
timestamp 0
transform 1 0 17572 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _0708_
timestamp 0
transform 1 0 19320 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0709_
timestamp 0
transform 1 0 26956 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0710_
timestamp 0
transform 1 0 26128 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0711_
timestamp 0
transform 1 0 26956 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0712_
timestamp 0
transform -1 0 26772 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0713_
timestamp 0
transform 1 0 22908 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0714_
timestamp 0
transform 1 0 21988 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0715_
timestamp 0
transform 1 0 19228 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0716_
timestamp 0
transform -1 0 18860 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0717_
timestamp 0
transform 1 0 21436 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0718_
timestamp 0
transform -1 0 21160 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0719_
timestamp 0
transform -1 0 27784 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0720_
timestamp 0
transform 1 0 28428 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0721_
timestamp 0
transform 1 0 26036 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0722_
timestamp 0
transform 1 0 26036 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0723_
timestamp 0
transform 1 0 26956 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0724_
timestamp 0
transform 1 0 26312 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0725_
timestamp 0
transform -1 0 18124 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _0726_
timestamp 0
transform 1 0 17296 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _0727_
timestamp 0
transform 1 0 19412 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0728_
timestamp 0
transform 1 0 29532 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0729_
timestamp 0
transform -1 0 28612 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0730_
timestamp 0
transform 1 0 29532 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0731_
timestamp 0
transform -1 0 29348 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0732_
timestamp 0
transform 1 0 24380 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0733_
timestamp 0
transform -1 0 23920 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0734_
timestamp 0
transform 1 0 20332 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0735_
timestamp 0
transform 1 0 20148 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0736_
timestamp 0
transform 1 0 26956 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0737_
timestamp 0
transform -1 0 26680 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0738_
timestamp 0
transform -1 0 30360 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0739_
timestamp 0
transform 1 0 30636 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0740_
timestamp 0
transform -1 0 29440 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0741_
timestamp 0
transform -1 0 30268 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0742_
timestamp 0
transform -1 0 29440 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0743_
timestamp 0
transform 1 0 31004 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0744_
timestamp 0
transform -1 0 14720 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _0745_
timestamp 0
transform -1 0 13984 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0746_
timestamp 0
transform 1 0 14076 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0747_
timestamp 0
transform -1 0 12512 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0748_
timestamp 0
transform 1 0 14628 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0749_
timestamp 0
transform -1 0 14076 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0750_
timestamp 0
transform 1 0 10120 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0751_
timestamp 0
transform -1 0 10764 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0752_
timestamp 0
transform 1 0 9476 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0753_
timestamp 0
transform -1 0 9016 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0754_
timestamp 0
transform -1 0 13984 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0755_
timestamp 0
transform -1 0 14352 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0756_
timestamp 0
transform 1 0 8832 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0757_
timestamp 0
transform -1 0 8832 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0758_
timestamp 0
transform 1 0 9476 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0759_
timestamp 0
transform 1 0 9200 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0760_
timestamp 0
transform 1 0 8924 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0761_
timestamp 0
transform -1 0 8464 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0762_
timestamp 0
transform -1 0 16560 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  _0763_
timestamp 0
transform 1 0 14720 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _0764_
timestamp 0
transform 1 0 15272 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0765_
timestamp 0
transform -1 0 16376 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0766_
timestamp 0
transform 1 0 16284 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0767_
timestamp 0
transform 1 0 14168 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0768_
timestamp 0
transform -1 0 13984 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0769_
timestamp 0
transform 1 0 7912 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0770_
timestamp 0
transform 1 0 7452 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0771_
timestamp 0
transform 1 0 8924 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0772_
timestamp 0
transform 1 0 8464 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0773_
timestamp 0
transform 1 0 15088 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0774_
timestamp 0
transform -1 0 14720 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0775_
timestamp 0
transform 1 0 7820 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0776_
timestamp 0
transform 1 0 7452 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0777_
timestamp 0
transform 1 0 8004 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0778_
timestamp 0
transform 1 0 7728 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0779_
timestamp 0
transform 1 0 8004 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0780_
timestamp 0
transform 1 0 7268 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0781_
timestamp 0
transform 1 0 16652 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__buf_4  _0782_
timestamp 0
transform 1 0 18032 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0783_
timestamp 0
transform 1 0 19228 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0784_
timestamp 0
transform -1 0 18400 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0785_
timestamp 0
transform 1 0 26956 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0786_
timestamp 0
transform -1 0 26036 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0787_
timestamp 0
transform 1 0 21896 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0788_
timestamp 0
transform -1 0 21712 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0789_
timestamp 0
transform 1 0 18124 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0790_
timestamp 0
transform -1 0 16560 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0791_
timestamp 0
transform 1 0 19596 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0792_
timestamp 0
transform 1 0 18216 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0793_
timestamp 0
transform -1 0 25300 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0794_
timestamp 0
transform 1 0 25852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0795_
timestamp 0
transform -1 0 28060 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0796_
timestamp 0
transform 1 0 28520 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0797_
timestamp 0
transform 1 0 26956 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0798_
timestamp 0
transform 1 0 26220 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _0799_
timestamp 0
transform 1 0 16836 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  _0800_
timestamp 0
transform 1 0 18860 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0801_
timestamp 0
transform 1 0 28612 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0802_
timestamp 0
transform -1 0 27968 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0803_
timestamp 0
transform -1 0 28796 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0804_
timestamp 0
transform -1 0 29256 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0805_
timestamp 0
transform 1 0 24380 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0806_
timestamp 0
transform -1 0 23368 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0807_
timestamp 0
transform 1 0 19320 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0808_
timestamp 0
transform -1 0 18860 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0809_
timestamp 0
transform 1 0 25944 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0810_
timestamp 0
transform 1 0 25760 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0811_
timestamp 0
transform -1 0 28888 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0812_
timestamp 0
transform 1 0 31096 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0813_
timestamp 0
transform 1 0 29164 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0814_
timestamp 0
transform -1 0 28612 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0815_
timestamp 0
transform -1 0 29992 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0816_
timestamp 0
transform 1 0 30728 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0817_
timestamp 0
transform -1 0 14720 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__buf_4  _0818_
timestamp 0
transform -1 0 13984 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0819_
timestamp 0
transform 1 0 13892 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0820_
timestamp 0
transform 1 0 13524 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0821_
timestamp 0
transform 1 0 14076 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0822_
timestamp 0
transform 1 0 13156 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0823_
timestamp 0
transform 1 0 7636 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0824_
timestamp 0
transform -1 0 7360 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0825_
timestamp 0
transform -1 0 9292 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0826_
timestamp 0
transform 1 0 9660 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0827_
timestamp 0
transform 1 0 12144 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0828_
timestamp 0
transform 1 0 12052 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0829_
timestamp 0
transform 1 0 7544 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0830_
timestamp 0
transform 1 0 6992 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0831_
timestamp 0
transform 1 0 7820 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0832_
timestamp 0
transform 1 0 7268 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0833_
timestamp 0
transform 1 0 7820 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0834_
timestamp 0
transform 1 0 7268 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0835_
timestamp 0
transform 1 0 16928 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  _0836_
timestamp 0
transform 1 0 18032 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _0837_
timestamp 0
transform 1 0 19228 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0838_
timestamp 0
transform 1 0 24472 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0839_
timestamp 0
transform -1 0 24288 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0840_
timestamp 0
transform 1 0 25668 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0841_
timestamp 0
transform 1 0 25576 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0842_
timestamp 0
transform 1 0 21896 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0843_
timestamp 0
transform -1 0 21436 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0844_
timestamp 0
transform 1 0 19228 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0845_
timestamp 0
transform 1 0 18032 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0846_
timestamp 0
transform 1 0 21160 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0847_
timestamp 0
transform 1 0 20976 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0848_
timestamp 0
transform -1 0 26220 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0849_
timestamp 0
transform -1 0 26588 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0850_
timestamp 0
transform 1 0 24380 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0851_
timestamp 0
transform -1 0 23920 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0852_
timestamp 0
transform 1 0 25116 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0853_
timestamp 0
transform 1 0 24012 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0854_
timestamp 0
transform 1 0 17388 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _0855_
timestamp 0
transform 1 0 19780 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0856_
timestamp 0
transform -1 0 21528 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0857_
timestamp 0
transform 1 0 21804 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0858_
timestamp 0
transform 1 0 25116 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0859_
timestamp 0
transform -1 0 24196 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0860_
timestamp 0
transform 1 0 21252 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0861_
timestamp 0
transform 1 0 21344 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0862_
timestamp 0
transform 1 0 18308 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0863_
timestamp 0
transform 1 0 17848 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0864_
timestamp 0
transform 1 0 19228 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0865_
timestamp 0
transform -1 0 19136 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0866_
timestamp 0
transform 1 0 22172 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0867_
timestamp 0
transform -1 0 21712 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0868_
timestamp 0
transform 1 0 23460 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0869_
timestamp 0
transform 1 0 23276 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0870_
timestamp 0
transform 1 0 24380 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0871_
timestamp 0
transform 1 0 23460 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _0872_
timestamp 0
transform -1 0 15272 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  _0873_
timestamp 0
transform -1 0 13432 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0874_
timestamp 0
transform 1 0 11500 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0875_
timestamp 0
transform 1 0 10948 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0876_
timestamp 0
transform 1 0 11960 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0877_
timestamp 0
transform 1 0 11684 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0878_
timestamp 0
transform 1 0 6164 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0879_
timestamp 0
transform -1 0 5980 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0880_
timestamp 0
transform 1 0 7176 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0881_
timestamp 0
transform -1 0 6256 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0882_
timestamp 0
transform 1 0 10856 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0883_
timestamp 0
transform 1 0 10580 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0884_
timestamp 0
transform 1 0 6348 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0885_
timestamp 0
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0886_
timestamp 0
transform -1 0 7176 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0887_
timestamp 0
transform 1 0 7544 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0888_
timestamp 0
transform 1 0 6624 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0889_
timestamp 0
transform -1 0 6256 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0890_
timestamp 0
transform -1 0 14076 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _0891_
timestamp 0
transform -1 0 8280 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0892_
timestamp 0
transform 1 0 3036 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0893_
timestamp 0
transform 1 0 2668 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0894_
timestamp 0
transform -1 0 7360 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0895_
timestamp 0
transform 1 0 6808 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0896_
timestamp 0
transform 1 0 3772 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0897_
timestamp 0
transform 1 0 2852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0898_
timestamp 0
transform 1 0 3772 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0899_
timestamp 0
transform -1 0 2208 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0900_
timestamp 0
transform 1 0 3772 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0901_
timestamp 0
transform -1 0 3036 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0902_
timestamp 0
transform 1 0 4232 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0903_
timestamp 0
transform -1 0 3680 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0904_
timestamp 0
transform 1 0 5428 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0905_
timestamp 0
transform 1 0 4324 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0906_
timestamp 0
transform 1 0 5244 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0907_
timestamp 0
transform 1 0 3956 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _0908_
timestamp 0
transform 1 0 16100 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  _0909_
timestamp 0
transform 1 0 18216 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0910_
timestamp 0
transform -1 0 17848 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0911_
timestamp 0
transform -1 0 18676 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0912_
timestamp 0
transform 1 0 24380 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0913_
timestamp 0
transform 1 0 23920 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0914_
timestamp 0
transform 1 0 20148 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0915_
timestamp 0
transform -1 0 19872 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0916_
timestamp 0
transform 1 0 17204 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0917_
timestamp 0
transform 1 0 17112 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0918_
timestamp 0
transform 1 0 17572 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0919_
timestamp 0
transform 1 0 17480 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0920_
timestamp 0
transform 1 0 22448 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0921_
timestamp 0
transform 1 0 22264 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0922_
timestamp 0
transform 1 0 23276 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0923_
timestamp 0
transform 1 0 23184 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0924_
timestamp 0
transform 1 0 24564 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0925_
timestamp 0
transform 1 0 23460 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0926_
timestamp 0
transform -1 0 15916 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _0927_
timestamp 0
transform -1 0 7636 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0928_
timestamp 0
transform 1 0 3772 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0929_
timestamp 0
transform 1 0 3772 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0930_
timestamp 0
transform -1 0 6808 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0931_
timestamp 0
transform 1 0 6992 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0932_
timestamp 0
transform 1 0 3956 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0933_
timestamp 0
transform 1 0 2576 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0934_
timestamp 0
transform -1 0 4876 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0935_
timestamp 0
transform 1 0 4968 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0936_
timestamp 0
transform 1 0 3772 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0937_
timestamp 0
transform 1 0 3036 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0938_
timestamp 0
transform 1 0 4876 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0939_
timestamp 0
transform -1 0 3404 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0940_
timestamp 0
transform -1 0 5428 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0941_
timestamp 0
transform 1 0 5336 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0942_
timestamp 0
transform 1 0 5060 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0943_
timestamp 0
transform -1 0 3588 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _0944_
timestamp 0
transform 1 0 15824 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  _0945_
timestamp 0
transform 1 0 18768 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0946_
timestamp 0
transform 1 0 17848 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0947_
timestamp 0
transform 1 0 17572 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0948_
timestamp 0
transform -1 0 27876 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0949_
timestamp 0
transform -1 0 28796 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0950_
timestamp 0
transform 1 0 20056 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0951_
timestamp 0
transform -1 0 19780 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0952_
timestamp 0
transform 1 0 16928 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0953_
timestamp 0
transform -1 0 16284 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0954_
timestamp 0
transform 1 0 18768 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0955_
timestamp 0
transform -1 0 17296 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0956_
timestamp 0
transform -1 0 24288 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0957_
timestamp 0
transform -1 0 24104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0958_
timestamp 0
transform 1 0 26956 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0959_
timestamp 0
transform 1 0 26404 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0960_
timestamp 0
transform 1 0 28428 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0961_
timestamp 0
transform 1 0 28152 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0962_
timestamp 0
transform -1 0 14720 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__buf_4  _0963_
timestamp 0
transform -1 0 13432 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0964_
timestamp 0
transform 1 0 12696 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0965_
timestamp 0
transform 1 0 12420 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0966_
timestamp 0
transform 1 0 14076 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0967_
timestamp 0
transform 1 0 13340 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0968_
timestamp 0
transform 1 0 6716 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0969_
timestamp 0
transform 1 0 5612 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0970_
timestamp 0
transform 1 0 6348 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0971_
timestamp 0
transform 1 0 5796 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0972_
timestamp 0
transform 1 0 12972 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0973_
timestamp 0
transform 1 0 11868 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0974_
timestamp 0
transform 1 0 7176 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0975_
timestamp 0
transform 1 0 6900 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0976_
timestamp 0
transform 1 0 8740 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0977_
timestamp 0
transform -1 0 8740 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0978_
timestamp 0
transform 1 0 6348 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0979_
timestamp 0
transform 1 0 6164 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _0980_
timestamp 0
transform 1 0 10580 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0981_
timestamp 0
transform 1 0 15640 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0982_
timestamp 0
transform 1 0 12144 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0983_
timestamp 0
transform 1 0 9016 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0984_
timestamp 0
transform 1 0 8648 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0985_
timestamp 0
transform 1 0 15272 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0986_
timestamp 0
transform 1 0 10304 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0987_
timestamp 0
transform 1 0 12880 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0988_
timestamp 0
transform 1 0 8924 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0989_
timestamp 0
transform 1 0 10764 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0990_
timestamp 0
transform 1 0 13800 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0991_
timestamp 0
transform 1 0 18768 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0992_
timestamp 0
transform 1 0 18400 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0993_
timestamp 0
transform -1 0 21344 0 1 30464
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0994_
timestamp 0
transform 1 0 15456 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0995_
timestamp 0
transform 1 0 16928 0 1 21760
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _0996_
timestamp 0
transform 1 0 16652 0 -1 22848
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0997_
timestamp 0
transform 1 0 18124 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0998_
timestamp 0
transform 1 0 16284 0 1 22848
box -38 -48 2154 592
use sky130_fd_sc_hd__dfxtp_1  _0999_
timestamp 0
transform 1 0 14628 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1000_
timestamp 0
transform 1 0 13892 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1001_
timestamp 0
transform 1 0 11500 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1002_
timestamp 0
transform 1 0 9936 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1003_
timestamp 0
transform 1 0 14076 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1004_
timestamp 0
transform 1 0 9752 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1005_
timestamp 0
transform 1 0 10764 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1006_
timestamp 0
transform 1 0 9936 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1007_
timestamp 0
transform 1 0 25852 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1008_
timestamp 0
transform 1 0 26680 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1009_
timestamp 0
transform 1 0 21804 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1010_
timestamp 0
transform 1 0 19136 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1011_
timestamp 0
transform -1 0 23276 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1012_
timestamp 0
transform -1 0 28428 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1013_
timestamp 0
transform 1 0 25760 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1014_
timestamp 0
transform 1 0 26036 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1015_
timestamp 0
transform 1 0 28612 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1016_
timestamp 0
transform 1 0 29532 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1017_
timestamp 0
transform 1 0 24840 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1018_
timestamp 0
transform 1 0 19320 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1019_
timestamp 0
transform 1 0 26956 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1020_
timestamp 0
transform 1 0 29532 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1021_
timestamp 0
transform -1 0 30636 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1022_
timestamp 0
transform -1 0 30728 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1023_
timestamp 0
transform 1 0 12512 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1024_
timestamp 0
transform 1 0 14076 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1025_
timestamp 0
transform -1 0 11224 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1026_
timestamp 0
transform 1 0 9016 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1027_
timestamp 0
transform -1 0 14628 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1028_
timestamp 0
transform 1 0 8924 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1029_
timestamp 0
transform 1 0 9016 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1030_
timestamp 0
transform -1 0 8832 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1031_
timestamp 0
transform 1 0 15088 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1032_
timestamp 0
transform 1 0 14076 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1033_
timestamp 0
transform 1 0 6992 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1034_
timestamp 0
transform 1 0 7360 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1035_
timestamp 0
transform 1 0 14720 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1036_
timestamp 0
transform 1 0 6992 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1037_
timestamp 0
transform 1 0 7268 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1038_
timestamp 0
transform 1 0 6532 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1039_
timestamp 0
transform 1 0 18768 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1040_
timestamp 0
transform 1 0 26036 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1041_
timestamp 0
transform 1 0 21804 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1042_
timestamp 0
transform 1 0 16560 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1043_
timestamp 0
transform 1 0 17664 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1044_
timestamp 0
transform -1 0 25392 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1045_
timestamp 0
transform 1 0 25392 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1046_
timestamp 0
transform 1 0 25944 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1047_
timestamp 0
transform 1 0 27968 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1048_
timestamp 0
transform 1 0 28796 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1049_
timestamp 0
transform 1 0 23368 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1050_
timestamp 0
transform 1 0 18860 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1051_
timestamp 0
transform 1 0 25484 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1052_
timestamp 0
transform -1 0 30360 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1053_
timestamp 0
transform 1 0 29532 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1054_
timestamp 0
transform -1 0 31004 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1055_
timestamp 0
transform -1 0 13892 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1056_
timestamp 0
transform 1 0 12788 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1057_
timestamp 0
transform 1 0 7084 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1058_
timestamp 0
transform 1 0 7360 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1059_
timestamp 0
transform 1 0 11500 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1060_
timestamp 0
transform 1 0 6440 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1061_
timestamp 0
transform 1 0 6716 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1062_
timestamp 0
transform 1 0 6992 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1063_
timestamp 0
transform 1 0 24380 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1064_
timestamp 0
transform 1 0 25208 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1065_
timestamp 0
transform 1 0 21436 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1066_
timestamp 0
transform 1 0 17664 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1067_
timestamp 0
transform 1 0 20240 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1068_
timestamp 0
transform 1 0 26220 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1069_
timestamp 0
transform 1 0 24380 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1070_
timestamp 0
transform 1 0 23644 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1071_
timestamp 0
transform -1 0 21712 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1072_
timestamp 0
transform 1 0 24380 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1073_
timestamp 0
transform 1 0 20700 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1074_
timestamp 0
transform 1 0 17480 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1075_
timestamp 0
transform 1 0 19228 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1076_
timestamp 0
transform 1 0 21804 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1077_
timestamp 0
transform 1 0 22908 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1078_
timestamp 0
transform 1 0 22816 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1079_
timestamp 0
transform 1 0 10580 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1080_
timestamp 0
transform 1 0 11408 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1081_
timestamp 0
transform 1 0 6900 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1082_
timestamp 0
transform 1 0 6348 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1083_
timestamp 0
transform 1 0 9936 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1084_
timestamp 0
transform 1 0 4968 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1085_
timestamp 0
transform 1 0 5244 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1086_
timestamp 0
transform 1 0 6348 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1087_
timestamp 0
transform 1 0 2300 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1088_
timestamp 0
transform 1 0 6348 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1089_
timestamp 0
transform 1 0 2484 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1090_
timestamp 0
transform 1 0 2208 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1091_
timestamp 0
transform 1 0 3956 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1092_
timestamp 0
transform 1 0 3772 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1093_
timestamp 0
transform 1 0 3864 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1094_
timestamp 0
transform 1 0 3772 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1095_
timestamp 0
transform 1 0 18308 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1096_
timestamp 0
transform 1 0 23644 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1097_
timestamp 0
transform 1 0 19872 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1098_
timestamp 0
transform 1 0 16836 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1099_
timestamp 0
transform 1 0 17204 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1100_
timestamp 0
transform 1 0 21804 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1101_
timestamp 0
transform 1 0 22816 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1102_
timestamp 0
transform 1 0 23092 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1103_
timestamp 0
transform 1 0 2208 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1104_
timestamp 0
transform -1 0 6992 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1105_
timestamp 0
transform 1 0 2484 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1106_
timestamp 0
transform 1 0 2576 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1107_
timestamp 0
transform 1 0 2484 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1108_
timestamp 0
transform 1 0 3404 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1109_
timestamp 0
transform 1 0 3956 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1110_
timestamp 0
transform 1 0 3588 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1111_
timestamp 0
transform 1 0 17296 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1112_
timestamp 0
transform -1 0 28980 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1113_
timestamp 0
transform 1 0 19780 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1114_
timestamp 0
transform 1 0 16652 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1115_
timestamp 0
transform 1 0 17296 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1116_
timestamp 0
transform 1 0 24380 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1117_
timestamp 0
transform 1 0 26036 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1118_
timestamp 0
transform 1 0 27508 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1119_
timestamp 0
transform 1 0 12144 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1120_
timestamp 0
transform 1 0 13156 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1121_
timestamp 0
transform 1 0 5244 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1122_
timestamp 0
transform 1 0 5428 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1123_
timestamp 0
transform 1 0 11776 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1124_
timestamp 0
transform 1 0 6532 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1125_
timestamp 0
transform 1 0 8924 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1126_
timestamp 0
transform 1 0 4784 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 0
transform -1 0 18492 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_clk
timestamp 0
transform -1 0 9476 0 -1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_clk
timestamp 0
transform -1 0 9936 0 1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_clk
timestamp 0
transform -1 0 13892 0 -1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_clk
timestamp 0
transform 1 0 12972 0 1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_clk
timestamp 0
transform -1 0 8556 0 -1 20672
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_clk
timestamp 0
transform 1 0 7912 0 -1 21760
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_clk
timestamp 0
transform 1 0 12144 0 1 20672
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_clk
timestamp 0
transform 1 0 11776 0 1 21760
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_clk
timestamp 0
transform -1 0 21620 0 -1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_clk
timestamp 0
transform 1 0 20516 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_clk
timestamp 0
transform 1 0 25392 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_clk
timestamp 0
transform 1 0 25852 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_clk
timestamp 0
transform -1 0 20792 0 1 21760
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_clk
timestamp 0
transform -1 0 21620 0 -1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_clk
timestamp 0
transform 1 0 25668 0 1 21760
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_clk
timestamp 0
transform 1 0 25300 0 -1 21760
box -38 -48 1050 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_9
timestamp 0
transform 1 0 1932 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_21
timestamp 0
transform 1 0 3036 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 0
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 0
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_41
timestamp 0
transform 1 0 4876 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_49
timestamp 0
transform 1 0 5612 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 0
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 0
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 0
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 0
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 0
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 0
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_119
timestamp 0
transform 1 0 12052 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_131
timestamp 0
transform 1 0 13156 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_139
timestamp 0
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 0
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_153
timestamp 0
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 0
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_169
timestamp 0
transform 1 0 16652 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_177
timestamp 0
transform 1 0 17388 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_184
timestamp 0
transform 1 0 18032 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_197
timestamp 0
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_209
timestamp 0
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_221
timestamp 0
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_225
timestamp 0
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_237
timestamp 0
transform 1 0 22908 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_247
timestamp 0
transform 1 0 23828 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_251
timestamp 0
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_253
timestamp 0
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_265
timestamp 0
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_277
timestamp 0
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_281
timestamp 0
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_293
timestamp 0
transform 1 0 28060 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_301
timestamp 0
transform 1 0 28796 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_309
timestamp 0
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_321
timestamp 0
transform 1 0 30636 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 0
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 0
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 0
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 0
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 0
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 0
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 0
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 0
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_81
timestamp 0
transform 1 0 8556 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_85
timestamp 0
transform 1 0 8924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_106
timestamp 0
transform 1 0 10856 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_116
timestamp 0
transform 1 0 11776 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_128
timestamp 0
transform 1 0 12880 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_133
timestamp 0
transform 1 0 13340 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_139
timestamp 0
transform 1 0 13892 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_151
timestamp 0
transform 1 0 14996 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_163
timestamp 0
transform 1 0 16100 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 0
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_172
timestamp 0
transform 1 0 16928 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_184
timestamp 0
transform 1 0 18032 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_196
timestamp 0
transform 1 0 19136 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_208
timestamp 0
transform 1 0 20240 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_220
timestamp 0
transform 1 0 21344 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 0
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_237
timestamp 0
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_249
timestamp 0
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_261
timestamp 0
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_273
timestamp 0
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 0
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_281
timestamp 0
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_293
timestamp 0
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_305
timestamp 0
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_317
timestamp 0
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_329
timestamp 0
transform 1 0 31372 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 0
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 0
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 0
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 0
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 0
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 0
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 0
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 0
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 0
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_85
timestamp 0
transform 1 0 8924 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_150
timestamp 0
transform 1 0 14904 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_178
timestamp 0
transform 1 0 17480 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_190
timestamp 0
transform 1 0 18584 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 0
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_209
timestamp 0
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_221
timestamp 0
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_233
timestamp 0
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_245
timestamp 0
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 0
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_253
timestamp 0
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_265
timestamp 0
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_277
timestamp 0
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_289
timestamp 0
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_301
timestamp 0
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_307
timestamp 0
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_309
timestamp 0
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_321
timestamp 0
transform 1 0 30636 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_329
timestamp 0
transform 1 0 31372 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 0
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 0
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 0
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 0
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 0
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 0
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_57
timestamp 0
transform 1 0 6348 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 0
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 0
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_121
timestamp 0
transform 1 0 12236 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_133
timestamp 0
transform 1 0 13340 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_145
timestamp 0
transform 1 0 14444 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_165
timestamp 0
transform 1 0 16284 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 0
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 0
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 0
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 0
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 0
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 0
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 0
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_237
timestamp 0
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_249
timestamp 0
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_261
timestamp 0
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_273
timestamp 0
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp 0
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_281
timestamp 0
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_293
timestamp 0
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_305
timestamp 0
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_317
timestamp 0
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_329
timestamp 0
transform 1 0 31372 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 0
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 0
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 0
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 0
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 0
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 0
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_96
timestamp 0
transform 1 0 9936 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_110
timestamp 0
transform 1 0 11224 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_122
timestamp 0
transform 1 0 12328 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_130
timestamp 0
transform 1 0 13064 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_134
timestamp 0
transform 1 0 13432 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 0
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_153
timestamp 0
transform 1 0 15180 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_174
timestamp 0
transform 1 0 17112 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_185
timestamp 0
transform 1 0 18124 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_193
timestamp 0
transform 1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 0
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_209
timestamp 0
transform 1 0 20332 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_229
timestamp 0
transform 1 0 22172 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_241
timestamp 0
transform 1 0 23276 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_249
timestamp 0
transform 1 0 24012 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 0
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_265
timestamp 0
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_277
timestamp 0
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_289
timestamp 0
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_301
timestamp 0
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_307
timestamp 0
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_309
timestamp 0
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_321
timestamp 0
transform 1 0 30636 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_329
timestamp 0
transform 1 0 31372 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 0
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 0
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 0
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 0
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 0
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 0
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 0
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_69
timestamp 0
transform 1 0 7452 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_97
timestamp 0
transform 1 0 10028 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_109
timestamp 0
transform 1 0 11132 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 0
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_125
timestamp 0
transform 1 0 12604 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_143
timestamp 0
transform 1 0 14260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_155
timestamp 0
transform 1 0 15364 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 0
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_169
timestamp 0
transform 1 0 16652 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_173
timestamp 0
transform 1 0 17020 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_177
timestamp 0
transform 1 0 17388 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_194
timestamp 0
transform 1 0 18952 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_200
timestamp 0
transform 1 0 19504 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 0
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_225
timestamp 0
transform 1 0 21804 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_234
timestamp 0
transform 1 0 22632 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_246
timestamp 0
transform 1 0 23736 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_258
timestamp 0
transform 1 0 24840 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_270
timestamp 0
transform 1 0 25944 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_278
timestamp 0
transform 1 0 26680 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_281
timestamp 0
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_293
timestamp 0
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_305
timestamp 0
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_317
timestamp 0
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_329
timestamp 0
transform 1 0 31372 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 0
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 0
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 0
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 0
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 0
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_53
timestamp 0
transform 1 0 5980 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_64
timestamp 0
transform 1 0 6992 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_76
timestamp 0
transform 1 0 8096 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 0
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 0
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_109
timestamp 0
transform 1 0 11132 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_128
timestamp 0
transform 1 0 12880 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_158
timestamp 0
transform 1 0 15640 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_170
timestamp 0
transform 1 0 16744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_205
timestamp 0
transform 1 0 19964 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_216
timestamp 0
transform 1 0 20976 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_228
timestamp 0
transform 1 0 22080 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_240
timestamp 0
transform 1 0 23184 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 0
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_269
timestamp 0
transform 1 0 25852 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_281
timestamp 0
transform 1 0 26956 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_293
timestamp 0
transform 1 0 28060 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_305
timestamp 0
transform 1 0 29164 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_309
timestamp 0
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_321
timestamp 0
transform 1 0 30636 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_329
timestamp 0
transform 1 0 31372 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_7
timestamp 0
transform 1 0 1748 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_19
timestamp 0
transform 1 0 2852 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_31
timestamp 0
transform 1 0 3956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_43
timestamp 0
transform 1 0 5060 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_49
timestamp 0
transform 1 0 5612 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_88
timestamp 0
transform 1 0 9200 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_100
timestamp 0
transform 1 0 10304 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_113
timestamp 0
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_135
timestamp 0
transform 1 0 13524 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_141
timestamp 0
transform 1 0 14076 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_153
timestamp 0
transform 1 0 15180 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_165
timestamp 0
transform 1 0 16284 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_169
timestamp 0
transform 1 0 16652 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_192
timestamp 0
transform 1 0 18768 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_201
timestamp 0
transform 1 0 19596 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_213
timestamp 0
transform 1 0 20700 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_232
timestamp 0
transform 1 0 22448 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_244
timestamp 0
transform 1 0 23552 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_278
timestamp 0
transform 1 0 26680 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_281
timestamp 0
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_293
timestamp 0
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_305
timestamp 0
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_317
timestamp 0
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_329
timestamp 0
transform 1 0 31372 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 0
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 0
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 0
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 0
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_41
timestamp 0
transform 1 0 4876 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_79
timestamp 0
transform 1 0 8372 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 0
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_85
timestamp 0
transform 1 0 8924 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_100
timestamp 0
transform 1 0 10304 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_105
timestamp 0
transform 1 0 10764 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_117
timestamp 0
transform 1 0 11868 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_129
timestamp 0
transform 1 0 12972 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_138
timestamp 0
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_157
timestamp 0
transform 1 0 15548 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_165
timestamp 0
transform 1 0 16284 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_178
timestamp 0
transform 1 0 17480 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_190
timestamp 0
transform 1 0 18584 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 0
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_209
timestamp 0
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_221
timestamp 0
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_233
timestamp 0
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_245
timestamp 0
transform 1 0 23644 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 0
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_277
timestamp 0
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_289
timestamp 0
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_301
timestamp 0
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_307
timestamp 0
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_309
timestamp 0
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_321
timestamp 0
transform 1 0 30636 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_329
timestamp 0
transform 1 0 31372 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 0
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 0
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 0
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_39
timestamp 0
transform 1 0 4692 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_47
timestamp 0
transform 1 0 5428 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_52
timestamp 0
transform 1 0 5888 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_110
timestamp 0
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 0
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_125
timestamp 0
transform 1 0 12604 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_164
timestamp 0
transform 1 0 16192 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 0
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_181
timestamp 0
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_193
timestamp 0
transform 1 0 18860 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_199
timestamp 0
transform 1 0 19412 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_219
timestamp 0
transform 1 0 21252 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_241
timestamp 0
transform 1 0 23276 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_253
timestamp 0
transform 1 0 24380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_265
timestamp 0
transform 1 0 25484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_277
timestamp 0
transform 1 0 26588 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_301
timestamp 0
transform 1 0 28796 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_313
timestamp 0
transform 1 0 29900 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_325
timestamp 0
transform 1 0 31004 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 0
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 0
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 0
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 0
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_41
timestamp 0
transform 1 0 4876 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_78
timestamp 0
transform 1 0 8280 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_85
timestamp 0
transform 1 0 8924 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_110
timestamp 0
transform 1 0 11224 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_122
timestamp 0
transform 1 0 12328 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_130
timestamp 0
transform 1 0 13064 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_136
timestamp 0
transform 1 0 13616 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_158
timestamp 0
transform 1 0 15640 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_166
timestamp 0
transform 1 0 16376 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_184
timestamp 0
transform 1 0 18032 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_197
timestamp 0
transform 1 0 19228 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_205
timestamp 0
transform 1 0 19964 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_223
timestamp 0
transform 1 0 21620 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_235
timestamp 0
transform 1 0 22724 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_244
timestamp 0
transform 1 0 23552 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_253
timestamp 0
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_265
timestamp 0
transform 1 0 25484 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_303
timestamp 0
transform 1 0 28980 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_307
timestamp 0
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_309
timestamp 0
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_321
timestamp 0
transform 1 0 30636 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 0
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 0
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 0
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 0
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_54
timestamp 0
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_57
timestamp 0
transform 1 0 6348 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_61
timestamp 0
transform 1 0 6716 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_70
timestamp 0
transform 1 0 7544 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_83
timestamp 0
transform 1 0 8740 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_87
timestamp 0
transform 1 0 9108 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_96
timestamp 0
transform 1 0 9936 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_107
timestamp 0
transform 1 0 10948 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 0
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 0
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_125
timestamp 0
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_137
timestamp 0
transform 1 0 13708 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_154
timestamp 0
transform 1 0 15272 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_202
timestamp 0
transform 1 0 19688 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_214
timestamp 0
transform 1 0 20792 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_222
timestamp 0
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_225
timestamp 0
transform 1 0 21804 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_233
timestamp 0
transform 1 0 22540 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_245
timestamp 0
transform 1 0 23644 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_257
timestamp 0
transform 1 0 24748 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_269
timestamp 0
transform 1 0 25852 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_281
timestamp 0
transform 1 0 26956 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_303
timestamp 0
transform 1 0 28980 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_315
timestamp 0
transform 1 0 30084 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_327
timestamp 0
transform 1 0 31188 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 0
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_15
timestamp 0
transform 1 0 2484 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_22
timestamp 0
transform 1 0 3128 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 0
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 0
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 0
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_65
timestamp 0
transform 1 0 7084 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_72
timestamp 0
transform 1 0 7728 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 0
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_97
timestamp 0
transform 1 0 10028 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_113
timestamp 0
transform 1 0 11500 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_126
timestamp 0
transform 1 0 12696 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_138
timestamp 0
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_141
timestamp 0
transform 1 0 14076 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_153
timestamp 0
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_165
timestamp 0
transform 1 0 16284 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_171
timestamp 0
transform 1 0 16836 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_197
timestamp 0
transform 1 0 19228 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_222
timestamp 0
transform 1 0 21528 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_230
timestamp 0
transform 1 0 22264 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_239
timestamp 0
transform 1 0 23092 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_243
timestamp 0
transform 1 0 23460 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_270
timestamp 0
transform 1 0 25944 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_274
timestamp 0
transform 1 0 26312 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_281
timestamp 0
transform 1 0 26956 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_293
timestamp 0
transform 1 0 28060 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_301
timestamp 0
transform 1 0 28796 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_306
timestamp 0
transform 1 0 29256 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_325
timestamp 0
transform 1 0 31004 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 0
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_31
timestamp 0
transform 1 0 3956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_43
timestamp 0
transform 1 0 5060 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 0
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_57
timestamp 0
transform 1 0 6348 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_63
timestamp 0
transform 1 0 6900 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_80
timestamp 0
transform 1 0 8464 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_92
timestamp 0
transform 1 0 9568 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_104
timestamp 0
transform 1 0 10672 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_108
timestamp 0
transform 1 0 11040 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_137
timestamp 0
transform 1 0 13708 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_169
timestamp 0
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_181
timestamp 0
transform 1 0 17756 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_189
timestamp 0
transform 1 0 18492 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_218
timestamp 0
transform 1 0 21160 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_225
timestamp 0
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_237
timestamp 0
transform 1 0 22908 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_274
timestamp 0
transform 1 0 26312 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_281
timestamp 0
transform 1 0 26956 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_289
timestamp 0
transform 1 0 27692 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_317
timestamp 0
transform 1 0 30268 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_327
timestamp 0
transform 1 0 31188 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 0
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_15
timestamp 0
transform 1 0 2484 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_19
timestamp 0
transform 1 0 2852 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 0
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_46
timestamp 0
transform 1 0 5336 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_58
timestamp 0
transform 1 0 6440 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_70
timestamp 0
transform 1 0 7544 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 0
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_93
timestamp 0
transform 1 0 9660 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_103
timestamp 0
transform 1 0 10580 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_110
timestamp 0
transform 1 0 11224 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_118
timestamp 0
transform 1 0 11960 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_130
timestamp 0
transform 1 0 13064 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_138
timestamp 0
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_150
timestamp 0
transform 1 0 14904 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_162
timestamp 0
transform 1 0 16008 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_174
timestamp 0
transform 1 0 17112 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_186
timestamp 0
transform 1 0 18216 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_194
timestamp 0
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_197
timestamp 0
transform 1 0 19228 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_223
timestamp 0
transform 1 0 21620 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_235
timestamp 0
transform 1 0 22724 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_243
timestamp 0
transform 1 0 23460 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_248
timestamp 0
transform 1 0 23920 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_270
timestamp 0
transform 1 0 25944 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_282
timestamp 0
transform 1 0 27048 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_294
timestamp 0
transform 1 0 28152 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_302
timestamp 0
transform 1 0 28888 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_307
timestamp 0
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_326
timestamp 0
transform 1 0 31096 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_330
timestamp 0
transform 1 0 31464 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 0
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 0
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_57
timestamp 0
transform 1 0 6348 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_68
timestamp 0
transform 1 0 7360 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_72
timestamp 0
transform 1 0 7728 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_94
timestamp 0
transform 1 0 9752 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_122
timestamp 0
transform 1 0 12328 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_139
timestamp 0
transform 1 0 13892 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_151
timestamp 0
transform 1 0 14996 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_163
timestamp 0
transform 1 0 16100 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_167
timestamp 0
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_169
timestamp 0
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_181
timestamp 0
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_193
timestamp 0
transform 1 0 18860 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_210
timestamp 0
transform 1 0 20424 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_222
timestamp 0
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_225
timestamp 0
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_237
timestamp 0
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_249
timestamp 0
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_261
timestamp 0
transform 1 0 25116 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_279
timestamp 0
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_290
timestamp 0
transform 1 0 27784 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_302
timestamp 0
transform 1 0 28888 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_314
timestamp 0
transform 1 0 29992 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_326
timestamp 0
transform 1 0 31096 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_330
timestamp 0
transform 1 0 31464 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_3
timestamp 0
transform 1 0 1380 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_46
timestamp 0
transform 1 0 5336 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_67
timestamp 0
transform 1 0 7268 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_107
timestamp 0
transform 1 0 10948 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_123
timestamp 0
transform 1 0 12420 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_168
timestamp 0
transform 1 0 16560 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_180
timestamp 0
transform 1 0 17664 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_187
timestamp 0
transform 1 0 18308 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_193
timestamp 0
transform 1 0 18860 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_221
timestamp 0
transform 1 0 21436 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_225
timestamp 0
transform 1 0 21804 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_242
timestamp 0
transform 1 0 23368 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_250
timestamp 0
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_253
timestamp 0
transform 1 0 24380 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_261
timestamp 0
transform 1 0 25116 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_302
timestamp 0
transform 1 0 28888 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_309
timestamp 0
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_321
timestamp 0
transform 1 0 30636 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_329
timestamp 0
transform 1 0 31372 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 0
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_15
timestamp 0
transform 1 0 2484 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_91
timestamp 0
transform 1 0 9476 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_103
timestamp 0
transform 1 0 10580 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 0
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_113
timestamp 0
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_125
timestamp 0
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_140
timestamp 0
transform 1 0 13984 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_169
timestamp 0
transform 1 0 16652 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_177
timestamp 0
transform 1 0 17388 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_223
timestamp 0
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_249
timestamp 0
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_261
timestamp 0
transform 1 0 25116 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_265
timestamp 0
transform 1 0 25484 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_269
timestamp 0
transform 1 0 25852 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_279
timestamp 0
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_289
timestamp 0
transform 1 0 27692 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_301
timestamp 0
transform 1 0 28796 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_313
timestamp 0
transform 1 0 29900 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_325
timestamp 0
transform 1 0 31004 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 0
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 0
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 0
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_29
timestamp 0
transform 1 0 3772 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_33
timestamp 0
transform 1 0 4140 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_45
timestamp 0
transform 1 0 5244 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_65
timestamp 0
transform 1 0 7084 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_76
timestamp 0
transform 1 0 8096 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 0
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_85
timestamp 0
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_99
timestamp 0
transform 1 0 10212 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_111
timestamp 0
transform 1 0 11316 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_123
timestamp 0
transform 1 0 12420 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_135
timestamp 0
transform 1 0 13524 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 0
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_141
timestamp 0
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_153
timestamp 0
transform 1 0 15180 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_174
timestamp 0
transform 1 0 17112 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_186
timestamp 0
transform 1 0 18216 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_194
timestamp 0
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_206
timestamp 0
transform 1 0 20056 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_215
timestamp 0
transform 1 0 20884 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_246
timestamp 0
transform 1 0 23736 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_253
timestamp 0
transform 1 0 24380 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_261
timestamp 0
transform 1 0 25116 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_275
timestamp 0
transform 1 0 26404 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_287
timestamp 0
transform 1 0 27508 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_299
timestamp 0
transform 1 0 28612 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_307
timestamp 0
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_318
timestamp 0
transform 1 0 30360 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_330
timestamp 0
transform 1 0 31464 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_9
timestamp 0
transform 1 0 1932 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_21
timestamp 0
transform 1 0 3036 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_33
timestamp 0
transform 1 0 4140 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_45
timestamp 0
transform 1 0 5244 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_53
timestamp 0
transform 1 0 5980 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_57
timestamp 0
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_69
timestamp 0
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_81
timestamp 0
transform 1 0 8556 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_105
timestamp 0
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 0
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_113
timestamp 0
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_125
timestamp 0
transform 1 0 12604 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_134
timestamp 0
transform 1 0 13432 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_144
timestamp 0
transform 1 0 14352 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_156
timestamp 0
transform 1 0 15456 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_169
timestamp 0
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_181
timestamp 0
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_193
timestamp 0
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_205
timestamp 0
transform 1 0 19964 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_222
timestamp 0
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_225
timestamp 0
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_230
timestamp 0
transform 1 0 22264 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_238
timestamp 0
transform 1 0 23000 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_249
timestamp 0
transform 1 0 24012 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_253
timestamp 0
transform 1 0 24380 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_263
timestamp 0
transform 1 0 25300 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_290
timestamp 0
transform 1 0 27784 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_323
timestamp 0
transform 1 0 30820 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 0
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 0
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 0
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_32
timestamp 0
transform 1 0 4048 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_44
timestamp 0
transform 1 0 5152 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_56
timestamp 0
transform 1 0 6256 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_68
timestamp 0
transform 1 0 7360 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_80
timestamp 0
transform 1 0 8464 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_85
timestamp 0
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_97
timestamp 0
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_109
timestamp 0
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_171
timestamp 0
transform 1 0 16836 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_183
timestamp 0
transform 1 0 17940 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_195
timestamp 0
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_205
timestamp 0
transform 1 0 19964 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_217
timestamp 0
transform 1 0 21068 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_229
timestamp 0
transform 1 0 22172 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_241
timestamp 0
transform 1 0 23276 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_285
timestamp 0
transform 1 0 27324 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_317
timestamp 0
transform 1 0 30268 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_329
timestamp 0
transform 1 0 31372 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_3
timestamp 0
transform 1 0 1380 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_11
timestamp 0
transform 1 0 2116 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_29
timestamp 0
transform 1 0 3772 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_46
timestamp 0
transform 1 0 5336 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_52
timestamp 0
transform 1 0 5888 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_57
timestamp 0
transform 1 0 6348 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_63
timestamp 0
transform 1 0 6900 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_67
timestamp 0
transform 1 0 7268 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_79
timestamp 0
transform 1 0 8372 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_91
timestamp 0
transform 1 0 9476 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_103
timestamp 0
transform 1 0 10580 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_110
timestamp 0
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_122
timestamp 0
transform 1 0 12328 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_148
timestamp 0
transform 1 0 14720 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_164
timestamp 0
transform 1 0 16192 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_173
timestamp 0
transform 1 0 17020 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_185
timestamp 0
transform 1 0 18124 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_210
timestamp 0
transform 1 0 20424 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_222
timestamp 0
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_231
timestamp 0
transform 1 0 22356 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_243
timestamp 0
transform 1 0 23460 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_255
timestamp 0
transform 1 0 24564 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_275
timestamp 0
transform 1 0 26404 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_279
timestamp 0
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_281
timestamp 0
transform 1 0 26956 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_293
timestamp 0
transform 1 0 28060 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_316
timestamp 0
transform 1 0 30176 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_320
timestamp 0
transform 1 0 30544 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_3
timestamp 0
transform 1 0 1380 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_11
timestamp 0
transform 1 0 2116 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_38
timestamp 0
transform 1 0 4600 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_82
timestamp 0
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_85
timestamp 0
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_97
timestamp 0
transform 1 0 10028 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_119
timestamp 0
transform 1 0 12052 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_138
timestamp 0
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_141
timestamp 0
transform 1 0 14076 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_171
timestamp 0
transform 1 0 16836 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_191
timestamp 0
transform 1 0 18676 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_195
timestamp 0
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_206
timestamp 0
transform 1 0 20056 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_224
timestamp 0
transform 1 0 21712 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_236
timestamp 0
transform 1 0 22816 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_248
timestamp 0
transform 1 0 23920 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_253
timestamp 0
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_265
timestamp 0
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_277
timestamp 0
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_289
timestamp 0
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_301
timestamp 0
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_307
timestamp 0
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_309
timestamp 0
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_321
timestamp 0
transform 1 0 30636 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_329
timestamp 0
transform 1 0 31372 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 0
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_15
timestamp 0
transform 1 0 2484 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_20
timestamp 0
transform 1 0 2944 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_38
timestamp 0
transform 1 0 4600 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_50
timestamp 0
transform 1 0 5704 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_66
timestamp 0
transform 1 0 7176 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_79
timestamp 0
transform 1 0 8372 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_83
timestamp 0
transform 1 0 8740 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_93
timestamp 0
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_105
timestamp 0
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 0
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_113
timestamp 0
transform 1 0 11500 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_119
timestamp 0
transform 1 0 12052 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_152
timestamp 0
transform 1 0 15088 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_164
timestamp 0
transform 1 0 16192 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_169
timestamp 0
transform 1 0 16652 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_175
timestamp 0
transform 1 0 17204 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_228
timestamp 0
transform 1 0 22080 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_238
timestamp 0
transform 1 0 23000 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_250
timestamp 0
transform 1 0 24104 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_262
timestamp 0
transform 1 0 25208 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_270
timestamp 0
transform 1 0 25944 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_297
timestamp 0
transform 1 0 28428 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_309
timestamp 0
transform 1 0 29532 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_321
timestamp 0
transform 1 0 30636 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_329
timestamp 0
transform 1 0 31372 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 0
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_15
timestamp 0
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 0
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_29
timestamp 0
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_41
timestamp 0
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_53
timestamp 0
transform 1 0 5980 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_59
timestamp 0
transform 1 0 6532 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_68
timestamp 0
transform 1 0 7360 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_79
timestamp 0
transform 1 0 8372 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_109
timestamp 0
transform 1 0 11132 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_117
timestamp 0
transform 1 0 11868 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_126
timestamp 0
transform 1 0 12696 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_138
timestamp 0
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_141
timestamp 0
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_153
timestamp 0
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_165
timestamp 0
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_177
timestamp 0
transform 1 0 17388 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_182
timestamp 0
transform 1 0 17848 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_191
timestamp 0
transform 1 0 18676 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_195
timestamp 0
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_205
timestamp 0
transform 1 0 19964 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_209
timestamp 0
transform 1 0 20332 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_217
timestamp 0
transform 1 0 21068 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_229
timestamp 0
transform 1 0 22172 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_249
timestamp 0
transform 1 0 24012 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_253
timestamp 0
transform 1 0 24380 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_261
timestamp 0
transform 1 0 25116 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_300
timestamp 0
transform 1 0 28704 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_309
timestamp 0
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_321
timestamp 0
transform 1 0 30636 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_329
timestamp 0
transform 1 0 31372 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 0
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_15
timestamp 0
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_27
timestamp 0
transform 1 0 3588 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_33
timestamp 0
transform 1 0 4140 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_43
timestamp 0
transform 1 0 5060 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp 0
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_57
timestamp 0
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_69
timestamp 0
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_81
timestamp 0
transform 1 0 8556 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_93
timestamp 0
transform 1 0 9660 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_111
timestamp 0
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_118
timestamp 0
transform 1 0 11960 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_130
timestamp 0
transform 1 0 13064 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_142
timestamp 0
transform 1 0 14168 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_150
timestamp 0
transform 1 0 14904 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_158
timestamp 0
transform 1 0 15640 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_166
timestamp 0
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_169
timestamp 0
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_181
timestamp 0
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_193
timestamp 0
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_205
timestamp 0
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_217
timestamp 0
transform 1 0 21068 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_264
timestamp 0
transform 1 0 25392 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_271
timestamp 0
transform 1 0 26036 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_277
timestamp 0
transform 1 0 26588 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_298
timestamp 0
transform 1 0 28520 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_310
timestamp 0
transform 1 0 29624 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_322
timestamp 0
transform 1 0 30728 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_330
timestamp 0
transform 1 0 31464 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 0
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_15
timestamp 0
transform 1 0 2484 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_21
timestamp 0
transform 1 0 3036 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_53
timestamp 0
transform 1 0 5980 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_61
timestamp 0
transform 1 0 6716 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_75
timestamp 0
transform 1 0 8004 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 0
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_85
timestamp 0
transform 1 0 8924 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_93
timestamp 0
transform 1 0 9660 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_118
timestamp 0
transform 1 0 11960 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_130
timestamp 0
transform 1 0 13064 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_138
timestamp 0
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_141
timestamp 0
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_153
timestamp 0
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_165
timestamp 0
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_177
timestamp 0
transform 1 0 17388 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_185
timestamp 0
transform 1 0 18124 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_189
timestamp 0
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_195
timestamp 0
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_197
timestamp 0
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_209
timestamp 0
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_221
timestamp 0
transform 1 0 21436 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_241
timestamp 0
transform 1 0 23276 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_272
timestamp 0
transform 1 0 26128 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_284
timestamp 0
transform 1 0 27232 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_296
timestamp 0
transform 1 0 28336 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_325
timestamp 0
transform 1 0 31004 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 0
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_15
timestamp 0
transform 1 0 2484 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_23
timestamp 0
transform 1 0 3220 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_50
timestamp 0
transform 1 0 5704 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_57
timestamp 0
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_89
timestamp 0
transform 1 0 9292 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_97
timestamp 0
transform 1 0 10028 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_102
timestamp 0
transform 1 0 10488 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_110
timestamp 0
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_113
timestamp 0
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_125
timestamp 0
transform 1 0 12604 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_129
timestamp 0
transform 1 0 12972 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_157
timestamp 0
transform 1 0 15548 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_166
timestamp 0
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_169
timestamp 0
transform 1 0 16652 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_177
timestamp 0
transform 1 0 17388 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_196
timestamp 0
transform 1 0 19136 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_208
timestamp 0
transform 1 0 20240 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_220
timestamp 0
transform 1 0 21344 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_225
timestamp 0
transform 1 0 21804 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_229
timestamp 0
transform 1 0 22172 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_233
timestamp 0
transform 1 0 22540 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_245
timestamp 0
transform 1 0 23644 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_250
timestamp 0
transform 1 0 24104 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_278
timestamp 0
transform 1 0 26680 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_281
timestamp 0
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_329
timestamp 0
transform 1 0 31372 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 0
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_15
timestamp 0
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 0
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_29
timestamp 0
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_41
timestamp 0
transform 1 0 4876 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_58
timestamp 0
transform 1 0 6440 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_80
timestamp 0
transform 1 0 8464 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_85
timestamp 0
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_97
timestamp 0
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_109
timestamp 0
transform 1 0 11132 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_117
timestamp 0
transform 1 0 11868 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_127
timestamp 0
transform 1 0 12788 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_144
timestamp 0
transform 1 0 14352 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_189
timestamp 0
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_195
timestamp 0
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_204
timestamp 0
transform 1 0 19872 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_217
timestamp 0
transform 1 0 21068 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_229
timestamp 0
transform 1 0 22172 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_241
timestamp 0
transform 1 0 23276 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_249
timestamp 0
transform 1 0 24012 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_261
timestamp 0
transform 1 0 25116 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_273
timestamp 0
transform 1 0 26220 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_285
timestamp 0
transform 1 0 27324 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_297
timestamp 0
transform 1 0 28428 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_318
timestamp 0
transform 1 0 30360 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_324
timestamp 0
transform 1 0 30912 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_330
timestamp 0
transform 1 0 31464 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_3
timestamp 0
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_15
timestamp 0
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_27
timestamp 0
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_39
timestamp 0
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_51
timestamp 0
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_55
timestamp 0
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_57
timestamp 0
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_72
timestamp 0
transform 1 0 7728 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_90
timestamp 0
transform 1 0 9384 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_102
timestamp 0
transform 1 0 10488 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_110
timestamp 0
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_113
timestamp 0
transform 1 0 11500 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_129
timestamp 0
transform 1 0 12972 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_147
timestamp 0
transform 1 0 14628 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_151
timestamp 0
transform 1 0 14996 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_161
timestamp 0
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_167
timestamp 0
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_169
timestamp 0
transform 1 0 16652 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_225
timestamp 0
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_237
timestamp 0
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_249
timestamp 0
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_261
timestamp 0
transform 1 0 25116 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_269
timestamp 0
transform 1 0 25852 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_279
timestamp 0
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_290
timestamp 0
transform 1 0 27784 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_299
timestamp 0
transform 1 0 28612 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_303
timestamp 0
transform 1 0 28980 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_308
timestamp 0
transform 1 0 29440 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_313
timestamp 0
transform 1 0 29900 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_325
timestamp 0
transform 1 0 31004 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_7
timestamp 0
transform 1 0 1748 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_15
timestamp 0
transform 1 0 2484 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_24
timestamp 0
transform 1 0 3312 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_53
timestamp 0
transform 1 0 5980 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_59
timestamp 0
transform 1 0 6532 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_77
timestamp 0
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_83
timestamp 0
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_85
timestamp 0
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_97
timestamp 0
transform 1 0 10028 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_115
timestamp 0
transform 1 0 11684 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_141
timestamp 0
transform 1 0 14076 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_176
timestamp 0
transform 1 0 17296 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_213
timestamp 0
transform 1 0 20700 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_242
timestamp 0
transform 1 0 23368 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_250
timestamp 0
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_253
timestamp 0
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_305
timestamp 0
transform 1 0 29164 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_309
timestamp 0
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_321
timestamp 0
transform 1 0 30636 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_329
timestamp 0
transform 1 0 31372 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_3
timestamp 0
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_47
timestamp 0
transform 1 0 5428 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_82
timestamp 0
transform 1 0 8648 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_94
timestamp 0
transform 1 0 9752 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_146
timestamp 0
transform 1 0 14536 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_155
timestamp 0
transform 1 0 15364 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_167
timestamp 0
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_169
timestamp 0
transform 1 0 16652 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_191
timestamp 0
transform 1 0 18676 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_196
timestamp 0
transform 1 0 19136 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_206
timestamp 0
transform 1 0 20056 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_241
timestamp 0
transform 1 0 23276 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_253
timestamp 0
transform 1 0 24380 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_265
timestamp 0
transform 1 0 25484 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_271
timestamp 0
transform 1 0 26036 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_278
timestamp 0
transform 1 0 26680 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_289
timestamp 0
transform 1 0 27692 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_301
timestamp 0
transform 1 0 28796 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_313
timestamp 0
transform 1 0 29900 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_325
timestamp 0
transform 1 0 31004 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_3
timestamp 0
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_15
timestamp 0
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 0
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_38
timestamp 0
transform 1 0 4600 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_48
timestamp 0
transform 1 0 5520 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_60
timestamp 0
transform 1 0 6624 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_80
timestamp 0
transform 1 0 8464 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_93
timestamp 0
transform 1 0 9660 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_105
timestamp 0
transform 1 0 10764 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_122
timestamp 0
transform 1 0 12328 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_126
timestamp 0
transform 1 0 12696 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_135
timestamp 0
transform 1 0 13524 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_139
timestamp 0
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_141
timestamp 0
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_153
timestamp 0
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_165
timestamp 0
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_177
timestamp 0
transform 1 0 17388 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_181
timestamp 0
transform 1 0 17756 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_195
timestamp 0
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_197
timestamp 0
transform 1 0 19228 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_205
timestamp 0
transform 1 0 19964 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_215
timestamp 0
transform 1 0 20884 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_219
timestamp 0
transform 1 0 21252 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_238
timestamp 0
transform 1 0 23000 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_246
timestamp 0
transform 1 0 23736 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_253
timestamp 0
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_265
timestamp 0
transform 1 0 25484 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_287
timestamp 0
transform 1 0 27508 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_295
timestamp 0
transform 1 0 28244 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_306
timestamp 0
transform 1 0 29256 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_309
timestamp 0
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_321
timestamp 0
transform 1 0 30636 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 0
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_15
timestamp 0
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_27
timestamp 0
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_39
timestamp 0
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_51
timestamp 0
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_55
timestamp 0
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_57
timestamp 0
transform 1 0 6348 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_65
timestamp 0
transform 1 0 7084 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_96
timestamp 0
transform 1 0 9936 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_108
timestamp 0
transform 1 0 11040 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_113
timestamp 0
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_125
timestamp 0
transform 1 0 12604 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_148
timestamp 0
transform 1 0 14720 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_160
timestamp 0
transform 1 0 15824 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_169
timestamp 0
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_181
timestamp 0
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_193
timestamp 0
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_205
timestamp 0
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_217
timestamp 0
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_223
timestamp 0
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_225
timestamp 0
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_237
timestamp 0
transform 1 0 22908 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_270
timestamp 0
transform 1 0 25944 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_277
timestamp 0
transform 1 0 26588 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_299
timestamp 0
transform 1 0 28612 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_305
timestamp 0
transform 1 0 29164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_322
timestamp 0
transform 1 0 30728 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_330
timestamp 0
transform 1 0 31464 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_3
timestamp 0
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_15
timestamp 0
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 0
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_29
timestamp 0
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_41
timestamp 0
transform 1 0 4876 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_58
timestamp 0
transform 1 0 6440 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_66
timestamp 0
transform 1 0 7176 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_94
timestamp 0
transform 1 0 9752 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_102
timestamp 0
transform 1 0 10488 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_112
timestamp 0
transform 1 0 11408 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_131
timestamp 0
transform 1 0 13156 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_139
timestamp 0
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_144
timestamp 0
transform 1 0 14352 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_156
timestamp 0
transform 1 0 15456 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_168
timestamp 0
transform 1 0 16560 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_180
timestamp 0
transform 1 0 17664 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_192
timestamp 0
transform 1 0 18768 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_197
timestamp 0
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_209
timestamp 0
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_221
timestamp 0
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_233
timestamp 0
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_245
timestamp 0
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_251
timestamp 0
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_253
timestamp 0
transform 1 0 24380 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_261
timestamp 0
transform 1 0 25116 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_278
timestamp 0
transform 1 0 26680 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_290
timestamp 0
transform 1 0 27784 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_328
timestamp 0
transform 1 0 31280 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_3
timestamp 0
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_15
timestamp 0
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_27
timestamp 0
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_39
timestamp 0
transform 1 0 4692 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_66
timestamp 0
transform 1 0 7176 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_93
timestamp 0
transform 1 0 9660 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_121
timestamp 0
transform 1 0 12236 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_135
timestamp 0
transform 1 0 13524 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_147
timestamp 0
transform 1 0 14628 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_159
timestamp 0
transform 1 0 15732 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_167
timestamp 0
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_169
timestamp 0
transform 1 0 16652 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_180
timestamp 0
transform 1 0 17664 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_192
timestamp 0
transform 1 0 18768 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_204
timestamp 0
transform 1 0 19872 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_216
timestamp 0
transform 1 0 20976 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_225
timestamp 0
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_237
timestamp 0
transform 1 0 22908 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_246
timestamp 0
transform 1 0 23736 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_274
timestamp 0
transform 1 0 26312 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_287
timestamp 0
transform 1 0 27508 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_299
timestamp 0
transform 1 0 28612 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_325
timestamp 0
transform 1 0 31004 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_3
timestamp 0
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_15
timestamp 0
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_27
timestamp 0
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_54
timestamp 0
transform 1 0 6072 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_58
timestamp 0
transform 1 0 6440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_76
timestamp 0
transform 1 0 8096 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_80
timestamp 0
transform 1 0 8464 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_85
timestamp 0
transform 1 0 8924 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_93
timestamp 0
transform 1 0 9660 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_109
timestamp 0
transform 1 0 11132 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_115
timestamp 0
transform 1 0 11684 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_127
timestamp 0
transform 1 0 12788 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_139
timestamp 0
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_141
timestamp 0
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_153
timestamp 0
transform 1 0 15180 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_161
timestamp 0
transform 1 0 15916 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_166
timestamp 0
transform 1 0 16376 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_195
timestamp 0
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_197
timestamp 0
transform 1 0 19228 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_214
timestamp 0
transform 1 0 20792 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_218
timestamp 0
transform 1 0 21160 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_224
timestamp 0
transform 1 0 21712 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_262
timestamp 0
transform 1 0 25208 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_266
timestamp 0
transform 1 0 25576 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_278
timestamp 0
transform 1 0 26680 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_290
timestamp 0
transform 1 0 27784 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_302
timestamp 0
transform 1 0 28888 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_317
timestamp 0
transform 1 0 30268 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_329
timestamp 0
transform 1 0 31372 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_3
timestamp 0
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_15
timestamp 0
transform 1 0 2484 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_23
timestamp 0
transform 1 0 3220 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_52
timestamp 0
transform 1 0 5888 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_57
timestamp 0
transform 1 0 6348 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_84
timestamp 0
transform 1 0 8832 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_96
timestamp 0
transform 1 0 9936 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_108
timestamp 0
transform 1 0 11040 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_113
timestamp 0
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_125
timestamp 0
transform 1 0 12604 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_138
timestamp 0
transform 1 0 13800 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_148
timestamp 0
transform 1 0 14720 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_156
timestamp 0
transform 1 0 15456 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_166
timestamp 0
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_195
timestamp 0
transform 1 0 19044 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_207
timestamp 0
transform 1 0 20148 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_223
timestamp 0
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_225
timestamp 0
transform 1 0 21804 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_229
timestamp 0
transform 1 0 22172 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_237
timestamp 0
transform 1 0 22908 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_264
timestamp 0
transform 1 0 25392 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_272
timestamp 0
transform 1 0 26128 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_281
timestamp 0
transform 1 0 26956 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_314
timestamp 0
transform 1 0 29992 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_326
timestamp 0
transform 1 0 31096 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_330
timestamp 0
transform 1 0 31464 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_3
timestamp 0
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_15
timestamp 0
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_27
timestamp 0
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_29
timestamp 0
transform 1 0 3772 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_34
timestamp 0
transform 1 0 4232 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_42
timestamp 0
transform 1 0 4968 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_60
timestamp 0
transform 1 0 6624 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_72
timestamp 0
transform 1 0 7728 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_93
timestamp 0
transform 1 0 9660 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_105
timestamp 0
transform 1 0 10764 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_117
timestamp 0
transform 1 0 11868 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_125
timestamp 0
transform 1 0 12604 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_138
timestamp 0
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_153
timestamp 0
transform 1 0 15180 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_161
timestamp 0
transform 1 0 15916 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_191
timestamp 0
transform 1 0 18676 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_197
timestamp 0
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_238
timestamp 0
transform 1 0 23000 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_242
timestamp 0
transform 1 0 23368 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_246
timestamp 0
transform 1 0 23736 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_253
timestamp 0
transform 1 0 24380 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_265
timestamp 0
transform 1 0 25484 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_269
timestamp 0
transform 1 0 25852 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_286
timestamp 0
transform 1 0 27416 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_303
timestamp 0
transform 1 0 28980 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_307
timestamp 0
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_309
timestamp 0
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_321
timestamp 0
transform 1 0 30636 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_329
timestamp 0
transform 1 0 31372 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_3
timestamp 0
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_15
timestamp 0
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_27
timestamp 0
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_39
timestamp 0
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_51
timestamp 0
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_55
timestamp 0
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_57
timestamp 0
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_69
timestamp 0
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_81
timestamp 0
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_93
timestamp 0
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_105
timestamp 0
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_111
timestamp 0
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_113
timestamp 0
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_125
timestamp 0
transform 1 0 12604 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_162
timestamp 0
transform 1 0 16008 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_169
timestamp 0
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_181
timestamp 0
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_193
timestamp 0
transform 1 0 18860 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_225
timestamp 0
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_237
timestamp 0
transform 1 0 22908 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_250
timestamp 0
transform 1 0 24104 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_260
timestamp 0
transform 1 0 25024 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_272
timestamp 0
transform 1 0 26128 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_276
timestamp 0
transform 1 0 26496 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_281
timestamp 0
transform 1 0 26956 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_285
timestamp 0
transform 1 0 27324 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_321
timestamp 0
transform 1 0 30636 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_329
timestamp 0
transform 1 0 31372 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_3
timestamp 0
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_15
timestamp 0
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_27
timestamp 0
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_29
timestamp 0
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_41
timestamp 0
transform 1 0 4876 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_47
timestamp 0
transform 1 0 5428 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_55
timestamp 0
transform 1 0 6164 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_67
timestamp 0
transform 1 0 7268 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_81
timestamp 0
transform 1 0 8556 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_85
timestamp 0
transform 1 0 8924 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_92
timestamp 0
transform 1 0 9568 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_102
timestamp 0
transform 1 0 10488 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_108
timestamp 0
transform 1 0 11040 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_121
timestamp 0
transform 1 0 12236 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_129
timestamp 0
transform 1 0 12972 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_139
timestamp 0
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_154
timestamp 0
transform 1 0 15272 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_162
timestamp 0
transform 1 0 16008 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_171
timestamp 0
transform 1 0 16836 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_183
timestamp 0
transform 1 0 17940 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_191
timestamp 0
transform 1 0 18676 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_195
timestamp 0
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_197
timestamp 0
transform 1 0 19228 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_214
timestamp 0
transform 1 0 20792 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_218
timestamp 0
transform 1 0 21160 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_226
timestamp 0
transform 1 0 21896 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_234
timestamp 0
transform 1 0 22632 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_247
timestamp 0
transform 1 0 23828 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_251
timestamp 0
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_253
timestamp 0
transform 1 0 24380 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_257
timestamp 0
transform 1 0 24748 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_262
timestamp 0
transform 1 0 25208 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_274
timestamp 0
transform 1 0 26312 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_286
timestamp 0
transform 1 0 27416 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_294
timestamp 0
transform 1 0 28152 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_325
timestamp 0
transform 1 0 31004 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_13
timestamp 0
transform 1 0 2300 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_25
timestamp 0
transform 1 0 3404 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_29
timestamp 0
transform 1 0 3772 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_49
timestamp 0
transform 1 0 5612 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_55
timestamp 0
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_57
timestamp 0
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_69
timestamp 0
transform 1 0 7452 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_84
timestamp 0
transform 1 0 8832 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_108
timestamp 0
transform 1 0 11040 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_122
timestamp 0
transform 1 0 12328 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_134
timestamp 0
transform 1 0 13432 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_141
timestamp 0
transform 1 0 14076 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_153
timestamp 0
transform 1 0 15180 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_165
timestamp 0
transform 1 0 16284 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_169
timestamp 0
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_181
timestamp 0
transform 1 0 17756 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_211
timestamp 0
transform 1 0 20516 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_223
timestamp 0
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_225
timestamp 0
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_237
timestamp 0
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_249
timestamp 0
transform 1 0 24012 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_258
timestamp 0
transform 1 0 24840 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_271
timestamp 0
transform 1 0 26036 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_279
timestamp 0
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_288
timestamp 0
transform 1 0 27600 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_296
timestamp 0
transform 1 0 28336 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_325
timestamp 0
transform 1 0 31004 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_3
timestamp 0
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_15
timestamp 0
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_27
timestamp 0
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_29
timestamp 0
transform 1 0 3772 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_64
timestamp 0
transform 1 0 6992 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_83
timestamp 0
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_100
timestamp 0
transform 1 0 10304 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_104
timestamp 0
transform 1 0 10672 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_129
timestamp 0
transform 1 0 12972 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_137
timestamp 0
transform 1 0 13708 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_141
timestamp 0
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_153
timestamp 0
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_165
timestamp 0
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_177
timestamp 0
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_189
timestamp 0
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_195
timestamp 0
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_200
timestamp 0
transform 1 0 19504 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_208
timestamp 0
transform 1 0 20240 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_214
timestamp 0
transform 1 0 20792 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_226
timestamp 0
transform 1 0 21896 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_238
timestamp 0
transform 1 0 23000 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_242
timestamp 0
transform 1 0 23368 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_262
timestamp 0
transform 1 0 25208 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_274
timestamp 0
transform 1 0 26312 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_286
timestamp 0
transform 1 0 27416 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_298
timestamp 0
transform 1 0 28520 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_306
timestamp 0
transform 1 0 29256 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_309
timestamp 0
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_321
timestamp 0
transform 1 0 30636 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_329
timestamp 0
transform 1 0 31372 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_3
timestamp 0
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_15
timestamp 0
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_27
timestamp 0
transform 1 0 3588 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_55
timestamp 0
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_66
timestamp 0
transform 1 0 7176 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_82
timestamp 0
transform 1 0 8648 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_90
timestamp 0
transform 1 0 9384 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_101
timestamp 0
transform 1 0 10396 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_109
timestamp 0
transform 1 0 11132 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_113
timestamp 0
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_125
timestamp 0
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_137
timestamp 0
transform 1 0 13708 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_160
timestamp 0
transform 1 0 15824 0 -1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_169
timestamp 0
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_181
timestamp 0
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_205
timestamp 0
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_217
timestamp 0
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_223
timestamp 0
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_225
timestamp 0
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_269
timestamp 0
transform 1 0 25852 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_289
timestamp 0
transform 1 0 27692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_301
timestamp 0
transform 1 0 28796 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_310
timestamp 0
transform 1 0 29624 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_322
timestamp 0
transform 1 0 30728 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_330
timestamp 0
transform 1 0 31464 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_3
timestamp 0
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_15
timestamp 0
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_27
timestamp 0
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_29
timestamp 0
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_41
timestamp 0
transform 1 0 4876 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_77
timestamp 0
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_83
timestamp 0
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_93
timestamp 0
transform 1 0 9660 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_105
timestamp 0
transform 1 0 10764 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_117
timestamp 0
transform 1 0 11868 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_125
timestamp 0
transform 1 0 12604 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_141
timestamp 0
transform 1 0 14076 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_145
timestamp 0
transform 1 0 14444 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_161
timestamp 0
transform 1 0 15916 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_169
timestamp 0
transform 1 0 16652 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_192
timestamp 0
transform 1 0 18768 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_209
timestamp 0
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_221
timestamp 0
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_233
timestamp 0
transform 1 0 22540 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_244
timestamp 0
transform 1 0 23552 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_248
timestamp 0
transform 1 0 23920 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_261
timestamp 0
transform 1 0 25116 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_267
timestamp 0
transform 1 0 25668 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_293
timestamp 0
transform 1 0 28060 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_305
timestamp 0
transform 1 0 29164 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_309
timestamp 0
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_321
timestamp 0
transform 1 0 30636 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_3
timestamp 0
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_15
timestamp 0
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_27
timestamp 0
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_39
timestamp 0
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_51
timestamp 0
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_55
timestamp 0
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_57
timestamp 0
transform 1 0 6348 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_69
timestamp 0
transform 1 0 7452 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_78
timestamp 0
transform 1 0 8280 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_86
timestamp 0
transform 1 0 9016 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_100
timestamp 0
transform 1 0 10304 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_113
timestamp 0
transform 1 0 11500 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_121
timestamp 0
transform 1 0 12236 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_147
timestamp 0
transform 1 0 14628 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_156
timestamp 0
transform 1 0 15456 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_204
timestamp 0
transform 1 0 19872 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_208
timestamp 0
transform 1 0 20240 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_216
timestamp 0
transform 1 0 20976 0 -1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_225
timestamp 0
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_237
timestamp 0
transform 1 0 22908 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_250
timestamp 0
transform 1 0 24104 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_262
timestamp 0
transform 1 0 25208 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_301
timestamp 0
transform 1 0 28796 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_313
timestamp 0
transform 1 0 29900 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_325
timestamp 0
transform 1 0 31004 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_3
timestamp 0
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_15
timestamp 0
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_27
timestamp 0
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_29
timestamp 0
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_41
timestamp 0
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_53
timestamp 0
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_71
timestamp 0
transform 1 0 7636 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_83
timestamp 0
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_85
timestamp 0
transform 1 0 8924 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_110
timestamp 0
transform 1 0 11224 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_122
timestamp 0
transform 1 0 12328 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_141
timestamp 0
transform 1 0 14076 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_145
timestamp 0
transform 1 0 14444 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_154
timestamp 0
transform 1 0 15272 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_162
timestamp 0
transform 1 0 16008 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_171
timestamp 0
transform 1 0 16836 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_195
timestamp 0
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_211
timestamp 0
transform 1 0 20516 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_221
timestamp 0
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_233
timestamp 0
transform 1 0 22540 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_261
timestamp 0
transform 1 0 25116 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_269
timestamp 0
transform 1 0 25852 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_295
timestamp 0
transform 1 0 28244 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_307
timestamp 0
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_309
timestamp 0
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_321
timestamp 0
transform 1 0 30636 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_329
timestamp 0
transform 1 0 31372 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_3
timestamp 0
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_15
timestamp 0
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_27
timestamp 0
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_39
timestamp 0
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_51
timestamp 0
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_55
timestamp 0
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_57
timestamp 0
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_69
timestamp 0
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_81
timestamp 0
transform 1 0 8556 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_92
timestamp 0
transform 1 0 9568 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_109
timestamp 0
transform 1 0 11132 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_113
timestamp 0
transform 1 0 11500 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_122
timestamp 0
transform 1 0 12328 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_152
timestamp 0
transform 1 0 15088 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_160
timestamp 0
transform 1 0 15824 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_178
timestamp 0
transform 1 0 17480 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_185
timestamp 0
transform 1 0 18124 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_197
timestamp 0
transform 1 0 19228 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_205
timestamp 0
transform 1 0 19964 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_214
timestamp 0
transform 1 0 20792 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_222
timestamp 0
transform 1 0 21528 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_225
timestamp 0
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_237
timestamp 0
transform 1 0 22908 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_243
timestamp 0
transform 1 0 23460 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_255
timestamp 0
transform 1 0 24564 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_267
timestamp 0
transform 1 0 25668 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_278
timestamp 0
transform 1 0 26680 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_281
timestamp 0
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_293
timestamp 0
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_305
timestamp 0
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_317
timestamp 0
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_329
timestamp 0
transform 1 0 31372 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_3
timestamp 0
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_15
timestamp 0
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_27
timestamp 0
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_29
timestamp 0
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_41
timestamp 0
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_53
timestamp 0
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_65
timestamp 0
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_77
timestamp 0
transform 1 0 8188 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_83
timestamp 0
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_101
timestamp 0
transform 1 0 10396 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_124
timestamp 0
transform 1 0 12512 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_136
timestamp 0
transform 1 0 13616 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_148
timestamp 0
transform 1 0 14720 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_160
timestamp 0
transform 1 0 15824 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_172
timestamp 0
transform 1 0 16928 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_184
timestamp 0
transform 1 0 18032 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_197
timestamp 0
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_209
timestamp 0
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_221
timestamp 0
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_233
timestamp 0
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_245
timestamp 0
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_251
timestamp 0
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_253
timestamp 0
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_265
timestamp 0
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_277
timestamp 0
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_289
timestamp 0
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_301
timestamp 0
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_307
timestamp 0
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_309
timestamp 0
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_321
timestamp 0
transform 1 0 30636 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_329
timestamp 0
transform 1 0 31372 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_3
timestamp 0
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_15
timestamp 0
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_27
timestamp 0
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_39
timestamp 0
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_51
timestamp 0
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_55
timestamp 0
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_57
timestamp 0
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_69
timestamp 0
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_81
timestamp 0
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_93
timestamp 0
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_105
timestamp 0
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_111
timestamp 0
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_113
timestamp 0
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_125
timestamp 0
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_137
timestamp 0
transform 1 0 13708 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_145
timestamp 0
transform 1 0 14444 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_150
timestamp 0
transform 1 0 14904 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_162
timestamp 0
transform 1 0 16008 0 -1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_169
timestamp 0
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_181
timestamp 0
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_193
timestamp 0
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_205
timestamp 0
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_217
timestamp 0
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_223
timestamp 0
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_225
timestamp 0
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_237
timestamp 0
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_249
timestamp 0
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_261
timestamp 0
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_273
timestamp 0
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_279
timestamp 0
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_281
timestamp 0
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_293
timestamp 0
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_305
timestamp 0
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_317
timestamp 0
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_329
timestamp 0
transform 1 0 31372 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_3
timestamp 0
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_15
timestamp 0
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_27
timestamp 0
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_29
timestamp 0
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_41
timestamp 0
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_53
timestamp 0
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_65
timestamp 0
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_77
timestamp 0
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_83
timestamp 0
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_85
timestamp 0
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_97
timestamp 0
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_109
timestamp 0
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_121
timestamp 0
transform 1 0 12236 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_146
timestamp 0
transform 1 0 14536 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_154
timestamp 0
transform 1 0 15272 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_160
timestamp 0
transform 1 0 15824 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_174
timestamp 0
transform 1 0 17112 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_183
timestamp 0
transform 1 0 17940 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_195
timestamp 0
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_197
timestamp 0
transform 1 0 19228 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_204
timestamp 0
transform 1 0 19872 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_216
timestamp 0
transform 1 0 20976 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_228
timestamp 0
transform 1 0 22080 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_240
timestamp 0
transform 1 0 23184 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_253
timestamp 0
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_265
timestamp 0
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_277
timestamp 0
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_289
timestamp 0
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_301
timestamp 0
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_307
timestamp 0
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_309
timestamp 0
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_321
timestamp 0
transform 1 0 30636 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_329
timestamp 0
transform 1 0 31372 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_3
timestamp 0
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_15
timestamp 0
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_27
timestamp 0
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_39
timestamp 0
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_51
timestamp 0
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_55
timestamp 0
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_57
timestamp 0
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_69
timestamp 0
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_81
timestamp 0
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_93
timestamp 0
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_105
timestamp 0
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_111
timestamp 0
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_113
timestamp 0
transform 1 0 11500 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_136
timestamp 0
transform 1 0 13616 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_142
timestamp 0
transform 1 0 14168 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_153
timestamp 0
transform 1 0 15180 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_157
timestamp 0
transform 1 0 15548 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_166
timestamp 0
transform 1 0 16376 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_187
timestamp 0
transform 1 0 18308 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_213
timestamp 0
transform 1 0 20700 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_221
timestamp 0
transform 1 0 21436 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_225
timestamp 0
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_237
timestamp 0
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_249
timestamp 0
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_261
timestamp 0
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_273
timestamp 0
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_279
timestamp 0
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_281
timestamp 0
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_293
timestamp 0
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_305
timestamp 0
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_317
timestamp 0
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_329
timestamp 0
transform 1 0 31372 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_7
timestamp 0
transform 1 0 1748 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_19
timestamp 0
transform 1 0 2852 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_27
timestamp 0
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_29
timestamp 0
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_41
timestamp 0
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_53
timestamp 0
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_65
timestamp 0
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_77
timestamp 0
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_83
timestamp 0
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_85
timestamp 0
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_97
timestamp 0
transform 1 0 10028 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_126
timestamp 0
transform 1 0 12696 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_130
timestamp 0
transform 1 0 13064 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_138
timestamp 0
transform 1 0 13800 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_144
timestamp 0
transform 1 0 14352 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_151
timestamp 0
transform 1 0 14996 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_155
timestamp 0
transform 1 0 15364 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_220
timestamp 0
transform 1 0 21344 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_232
timestamp 0
transform 1 0 22448 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_244
timestamp 0
transform 1 0 23552 0 1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_253
timestamp 0
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_265
timestamp 0
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_277
timestamp 0
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_289
timestamp 0
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_301
timestamp 0
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_307
timestamp 0
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_309
timestamp 0
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_321
timestamp 0
transform 1 0 30636 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_329
timestamp 0
transform 1 0 31372 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_3
timestamp 0
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_15
timestamp 0
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_27
timestamp 0
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_39
timestamp 0
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_51
timestamp 0
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_55
timestamp 0
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_57
timestamp 0
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_69
timestamp 0
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_81
timestamp 0
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_93
timestamp 0
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_105
timestamp 0
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_111
timestamp 0
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_113
timestamp 0
transform 1 0 11500 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_121
timestamp 0
transform 1 0 12236 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_133
timestamp 0
transform 1 0 13340 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_158
timestamp 0
transform 1 0 15640 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_166
timestamp 0
transform 1 0 16376 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_169
timestamp 0
transform 1 0 16652 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_185
timestamp 0
transform 1 0 18124 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_209
timestamp 0
transform 1 0 20332 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_221
timestamp 0
transform 1 0 21436 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_225
timestamp 0
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_237
timestamp 0
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_249
timestamp 0
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_261
timestamp 0
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_273
timestamp 0
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_279
timestamp 0
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_281
timestamp 0
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_293
timestamp 0
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_305
timestamp 0
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_317
timestamp 0
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_329
timestamp 0
transform 1 0 31372 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_3
timestamp 0
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_15
timestamp 0
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_27
timestamp 0
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_29
timestamp 0
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_41
timestamp 0
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_53
timestamp 0
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_65
timestamp 0
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_77
timestamp 0
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_83
timestamp 0
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_85
timestamp 0
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_97
timestamp 0
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_109
timestamp 0
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_121
timestamp 0
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_133
timestamp 0
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_139
timestamp 0
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_141
timestamp 0
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_153
timestamp 0
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_165
timestamp 0
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_177
timestamp 0
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_189
timestamp 0
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_195
timestamp 0
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_205
timestamp 0
transform 1 0 19964 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_217
timestamp 0
transform 1 0 21068 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_229
timestamp 0
transform 1 0 22172 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_241
timestamp 0
transform 1 0 23276 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_249
timestamp 0
transform 1 0 24012 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_253
timestamp 0
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_265
timestamp 0
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_277
timestamp 0
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_289
timestamp 0
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_301
timestamp 0
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_307
timestamp 0
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_309
timestamp 0
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_321
timestamp 0
transform 1 0 30636 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_329
timestamp 0
transform 1 0 31372 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_6
timestamp 0
transform 1 0 1656 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_18
timestamp 0
transform 1 0 2760 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_26
timestamp 0
transform 1 0 3496 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_29
timestamp 0
transform 1 0 3772 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_41
timestamp 0
transform 1 0 4876 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_53
timestamp 0
transform 1 0 5980 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_57
timestamp 0
transform 1 0 6348 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_65
timestamp 0
transform 1 0 7084 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_70
timestamp 0
transform 1 0 7544 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_82
timestamp 0
transform 1 0 8648 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_85
timestamp 0
transform 1 0 8924 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_97
timestamp 0
transform 1 0 10028 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_109
timestamp 0
transform 1 0 11132 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_113
timestamp 0
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_125
timestamp 0
transform 1 0 12604 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_133
timestamp 0
transform 1 0 13340 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_139
timestamp 0
transform 1 0 13892 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_141
timestamp 0
transform 1 0 14076 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_153
timestamp 0
transform 1 0 15180 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_165
timestamp 0
transform 1 0 16284 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_169
timestamp 0
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_181
timestamp 0
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_193
timestamp 0
transform 1 0 18860 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_203
timestamp 0
transform 1 0 19780 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_215
timestamp 0
transform 1 0 20884 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_223
timestamp 0
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_225
timestamp 0
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_237
timestamp 0
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_249
timestamp 0
transform 1 0 24012 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_253
timestamp 0
transform 1 0 24380 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_261
timestamp 0
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_273
timestamp 0
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_279
timestamp 0
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_281
timestamp 0
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_293
timestamp 0
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_305
timestamp 0
transform 1 0 29164 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_309
timestamp 0
transform 1 0 29532 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_317
timestamp 0
transform 1 0 30268 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_322
timestamp 0
transform 1 0 30728 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_330
timestamp 0
transform 1 0 31464 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp 0
transform -1 0 16836 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 0
transform -1 0 12972 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 0
transform -1 0 16008 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 0
transform -1 0 16100 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 0
transform -1 0 12236 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 0
transform -1 0 11960 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 0
transform -1 0 14076 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 0
transform -1 0 15640 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 0
transform -1 0 9384 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 0
transform 1 0 18400 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 0
transform -1 0 22724 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 0
transform -1 0 20884 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 0
transform 1 0 24564 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 0
transform -1 0 5336 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 0
transform -1 0 13708 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 0
transform -1 0 30268 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 0
transform -1 0 14352 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 0
transform 1 0 20976 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 0
transform 1 0 11684 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 0
transform -1 0 26036 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 0
transform -1 0 16928 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 0
transform -1 0 24012 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 0
transform -1 0 15088 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 0
transform -1 0 23644 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 0
transform -1 0 14536 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 0
transform -1 0 12052 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 0
transform -1 0 28612 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 0
transform -1 0 28520 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 0
transform -1 0 26128 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 0
transform -1 0 24012 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 0
transform -1 0 25944 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 0
transform -1 0 17112 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 0
transform -1 0 30820 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 0
transform -1 0 25116 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 0
transform 1 0 24748 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 0
transform -1 0 8740 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 0
transform -1 0 9660 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp 0
transform -1 0 19964 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 0
transform -1 0 30728 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp 0
transform -1 0 21528 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 0
transform -1 0 29440 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 0
transform -1 0 31096 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 0
transform -1 0 9660 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 0
transform -1 0 11224 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp 0
transform -1 0 5980 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp 0
transform -1 0 28428 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 0
transform -1 0 20884 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold48
timestamp 0
transform -1 0 30176 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp 0
transform -1 0 13524 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold50
timestamp 0
transform -1 0 19964 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp 0
transform 1 0 28428 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold52
timestamp 0
transform -1 0 27692 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp 0
transform -1 0 29164 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold54
timestamp 0
transform -1 0 23552 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold55
timestamp 0
transform -1 0 28520 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold56
timestamp 0
transform -1 0 21712 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold57
timestamp 0
transform -1 0 25944 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold58
timestamp 0
transform -1 0 28152 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold59
timestamp 0
transform -1 0 15640 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold60
timestamp 0
transform -1 0 20976 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold61
timestamp 0
transform -1 0 16284 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold62
timestamp 0
transform -1 0 24012 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold63
timestamp 0
transform -1 0 22632 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold64
timestamp 0
transform -1 0 28612 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold65
timestamp 0
transform -1 0 5980 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold66
timestamp 0
transform -1 0 5796 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold67
timestamp 0
transform -1 0 29992 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold68
timestamp 0
transform -1 0 20792 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold69
timestamp 0
transform -1 0 19044 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold70
timestamp 0
transform -1 0 28888 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold71
timestamp 0
transform -1 0 11132 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold72
timestamp 0
transform -1 0 8648 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold73
timestamp 0
transform -1 0 13524 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold74
timestamp 0
transform -1 0 21620 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold75
timestamp 0
transform -1 0 9660 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold76
timestamp 0
transform -1 0 31188 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold77
timestamp 0
transform -1 0 12696 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold78
timestamp 0
transform -1 0 9660 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold79
timestamp 0
transform -1 0 4692 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold80
timestamp 0
transform -1 0 28612 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold81
timestamp 0
transform -1 0 26036 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold82
timestamp 0
transform -1 0 4600 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold83
timestamp 0
transform -1 0 26680 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold84
timestamp 0
transform -1 0 21160 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold85
timestamp 0
transform -1 0 29992 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold86
timestamp 0
transform -1 0 18768 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold87
timestamp 0
transform -1 0 8188 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold88
timestamp 0
transform -1 0 9660 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold89
timestamp 0
transform -1 0 18492 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold90
timestamp 0
transform -1 0 27692 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold91
timestamp 0
transform -1 0 28244 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold92
timestamp 0
transform 1 0 8556 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold93
timestamp 0
transform 1 0 10120 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold94
timestamp 0
transform -1 0 8096 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold95
timestamp 0
transform -1 0 20884 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold96
timestamp 0
transform 1 0 24380 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold97
timestamp 0
transform -1 0 4968 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold98
timestamp 0
transform -1 0 23000 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold99
timestamp 0
transform -1 0 5520 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold100
timestamp 0
transform -1 0 6992 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold101
timestamp 0
transform -1 0 5336 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold102
timestamp 0
transform -1 0 25116 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold103
timestamp 0
transform -1 0 26036 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold104
timestamp 0
transform -1 0 10028 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold105
timestamp 0
transform -1 0 19688 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold106
timestamp 0
transform -1 0 7452 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold107
timestamp 0
transform -1 0 11224 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold108
timestamp 0
transform -1 0 25944 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold109
timestamp 0
transform -1 0 6164 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold110
timestamp 0
transform -1 0 7360 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold111
timestamp 0
transform -1 0 5520 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold112
timestamp 0
transform -1 0 28520 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold113
timestamp 0
transform -1 0 10672 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold114
timestamp 0
transform -1 0 15640 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold115
timestamp 0
transform -1 0 28060 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold116
timestamp 0
transform -1 0 31004 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold117
timestamp 0
transform 1 0 5520 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold118
timestamp 0
transform -1 0 8280 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold119
timestamp 0
transform -1 0 8740 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold120
timestamp 0
transform -1 0 5336 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold121
timestamp 0
transform -1 0 10488 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold122
timestamp 0
transform -1 0 6164 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold123
timestamp 0
transform -1 0 7268 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold124
timestamp 0
transform -1 0 19964 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold125
timestamp 0
transform -1 0 16192 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold126
timestamp 0
transform -1 0 9660 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold127
timestamp 0
transform -1 0 12328 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold128
timestamp 0
transform -1 0 8556 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold129
timestamp 0
transform -1 0 13064 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold130
timestamp 0
transform -1 0 7544 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold131
timestamp 0
transform -1 0 18124 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold132
timestamp 0
transform -1 0 12236 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold133
timestamp 0
transform -1 0 19964 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold134
timestamp 0
transform -1 0 19136 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold135
timestamp 0
transform -1 0 11224 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  input1
timestamp 0
transform 1 0 1380 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input2
timestamp 0
transform 1 0 29072 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input3
timestamp 0
transform 1 0 1380 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input4
timestamp 0
transform 1 0 1380 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input5
timestamp 0
transform 1 0 7176 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input6
timestamp 0
transform 1 0 12972 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input7
timestamp 0
transform 1 0 30360 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input8
timestamp 0
transform -1 0 31556 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input9
timestamp 0
transform 1 0 1380 0 -1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input10
timestamp 0
transform 1 0 1380 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input11
timestamp 0
transform -1 0 31556 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  max_cap1
timestamp 0
transform 1 0 23184 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  max_cap2
timestamp 0
transform 1 0 22908 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  max_cap23
timestamp 0
transform 1 0 14628 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output12
timestamp 0
transform 1 0 23276 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output13
timestamp 0
transform -1 0 1932 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output14
timestamp 0
transform -1 0 6256 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output15
timestamp 0
transform -1 0 1932 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output16
timestamp 0
transform 1 0 31188 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output17
timestamp 0
transform -1 0 12052 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output18
timestamp 0
transform 1 0 31188 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output19
timestamp 0
transform 1 0 31004 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output20
timestamp 0
transform 1 0 19228 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output21
timestamp 0
transform 1 0 24564 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output22
timestamp 0
transform 1 0 17480 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 0
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 0
transform -1 0 31832 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 0
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 0
transform -1 0 31832 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 0
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 0
transform -1 0 31832 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 0
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 0
transform -1 0 31832 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 0
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 0
transform -1 0 31832 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 0
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 0
transform -1 0 31832 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 0
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 0
transform -1 0 31832 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 0
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 0
transform -1 0 31832 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 0
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 0
transform -1 0 31832 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 0
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 0
transform -1 0 31832 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 0
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 0
transform -1 0 31832 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 0
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 0
transform -1 0 31832 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 0
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 0
transform -1 0 31832 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 0
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 0
transform -1 0 31832 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 0
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 0
transform -1 0 31832 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 0
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 0
transform -1 0 31832 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 0
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 0
transform -1 0 31832 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 0
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 0
transform -1 0 31832 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 0
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 0
transform -1 0 31832 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 0
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 0
transform -1 0 31832 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 0
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 0
transform -1 0 31832 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 0
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 0
transform -1 0 31832 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 0
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 0
transform -1 0 31832 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 0
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 0
transform -1 0 31832 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 0
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 0
transform -1 0 31832 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 0
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 0
transform -1 0 31832 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 0
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 0
transform -1 0 31832 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 0
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 0
transform -1 0 31832 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 0
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 0
transform -1 0 31832 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 0
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 0
transform -1 0 31832 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 0
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 0
transform -1 0 31832 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 0
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 0
transform -1 0 31832 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 0
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 0
transform -1 0 31832 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 0
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 0
transform -1 0 31832 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 0
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 0
transform -1 0 31832 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 0
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 0
transform -1 0 31832 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 0
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 0
transform -1 0 31832 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 0
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 0
transform -1 0 31832 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 0
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 0
transform -1 0 31832 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 0
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 0
transform -1 0 31832 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 0
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 0
transform -1 0 31832 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 0
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 0
transform -1 0 31832 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 0
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 0
transform -1 0 31832 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 0
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 0
transform -1 0 31832 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 0
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 0
transform -1 0 31832 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 0
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 0
transform -1 0 31832 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 0
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 0
transform -1 0 31832 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 0
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 0
transform -1 0 31832 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 0
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 0
transform -1 0 31832 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 0
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 0
transform -1 0 31832 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 0
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 0
transform -1 0 31832 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 0
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 0
transform -1 0 31832 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 0
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 0
transform -1 0 31832 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 0
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 0
transform -1 0 31832 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 0
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 0
transform -1 0 31832 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 0
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 0
transform -1 0 31832 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 0
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 0
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 0
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 0
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 0
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 0
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 0
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 0
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 0
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 0
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 0
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 0
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 0
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 0
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 0
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 0
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 0
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 0
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 0
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 0
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 0
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 0
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 0
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 0
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 0
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 0
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 0
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 0
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 0
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 0
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 0
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 0
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 0
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 0
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 0
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 0
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 0
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 0
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 0
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 0
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 0
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 0
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 0
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 0
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 0
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 0
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 0
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 0
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 0
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 0
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 0
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 0
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 0
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 0
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 0
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 0
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 0
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 0
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 0
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 0
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 0
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 0
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 0
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 0
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 0
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 0
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 0
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 0
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 0
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 0
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 0
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 0
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 0
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 0
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 0
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 0
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 0
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 0
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 0
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 0
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 0
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 0
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 0
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 0
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 0
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 0
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 0
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 0
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 0
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 0
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 0
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 0
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 0
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 0
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 0
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 0
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 0
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 0
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 0
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 0
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 0
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 0
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 0
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 0
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 0
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 0
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 0
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 0
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 0
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 0
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 0
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 0
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 0
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 0
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 0
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 0
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 0
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 0
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 0
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 0
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 0
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 0
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 0
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 0
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 0
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 0
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 0
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 0
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 0
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 0
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 0
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 0
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 0
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 0
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 0
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 0
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 0
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 0
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 0
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 0
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 0
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 0
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 0
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 0
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 0
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 0
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 0
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 0
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 0
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 0
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 0
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 0
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 0
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 0
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 0
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 0
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 0
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 0
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 0
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 0
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 0
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 0
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 0
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 0
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 0
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 0
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 0
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 0
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 0
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 0
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 0
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 0
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 0
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 0
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 0
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 0
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 0
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 0
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 0
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 0
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 0
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 0
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 0
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 0
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 0
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 0
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 0
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 0
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 0
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 0
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 0
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 0
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 0
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 0
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 0
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 0
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 0
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 0
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 0
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 0
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 0
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 0
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 0
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 0
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 0
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 0
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 0
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 0
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 0
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 0
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 0
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 0
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 0
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 0
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 0
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 0
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 0
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 0
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 0
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 0
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 0
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 0
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 0
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 0
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 0
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 0
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 0
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 0
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 0
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 0
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 0
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 0
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 0
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 0
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 0
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 0
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 0
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 0
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 0
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 0
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 0
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 0
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 0
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 0
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 0
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 0
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 0
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 0
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 0
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 0
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 0
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 0
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 0
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 0
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 0
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 0
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 0
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 0
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 0
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 0
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 0
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 0
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 0
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 0
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 0
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 0
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 0
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 0
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 0
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 0
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 0
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 0
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 0
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 0
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 0
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 0
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 0
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 0
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 0
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 0
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 0
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 0
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 0
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 0
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 0
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 0
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 0
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 0
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 0
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 0
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 0
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 0
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 0
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 0
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 0
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 0
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 0
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 0
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 0
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 0
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 0
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 0
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 0
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 0
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 0
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 0
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 0
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 0
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 0
transform 1 0 3680 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 0
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 0
transform 1 0 8832 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 0
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 0
transform 1 0 13984 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 0
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 0
transform 1 0 19136 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 0
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 0
transform 1 0 24288 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 0
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 0
transform 1 0 29440 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  wire3
timestamp 0
transform 1 0 26956 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  wire4
timestamp 0
transform 1 0 27508 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  wire24
timestamp 0
transform 1 0 24656 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  wire25
timestamp 0
transform 1 0 24840 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  wire26
timestamp 0
transform 1 0 29072 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  wire27
timestamp 0
transform 1 0 29532 0 -1 18496
box -38 -48 406 592
<< labels >>
rlabel metal1 s 16468 32640 16468 32640 4 VGND
rlabel metal2 s 16468 32096 16468 32096 4 VPWR
rlabel metal1 s 13938 30906 13938 30906 4 _0000_
rlabel metal1 s 12266 28458 12266 28458 4 _0001_
rlabel metal1 s 16744 3162 16744 3162 4 _0002_
rlabel metal2 s 13754 3298 13754 3298 4 _0003_
rlabel metal2 s 9890 3230 9890 3230 4 _0004_
rlabel metal1 s 10403 12886 10403 12886 4 _0005_
rlabel metal1 s 16468 3162 16468 3162 4 _0006_
rlabel metal2 s 11638 3298 11638 3298 4 _0007_
rlabel metal2 s 14214 20638 14214 20638 4 _0008_
rlabel metal1 s 10633 24786 10633 24786 4 _0009_
rlabel metal1 s 12190 30743 12190 30743 4 _0010_
rlabel metal2 s 14858 31144 14858 31144 4 _0011_
rlabel metal2 s 19734 30056 19734 30056 4 _0012_
rlabel metal2 s 19458 30600 19458 30600 4 _0013_
rlabel metal1 s 18768 30022 18768 30022 4 _0014_
rlabel metal2 s 16882 30906 16882 30906 4 _0015_
rlabel metal1 s 18453 21998 18453 21998 4 _0016_
rlabel metal1 s 18545 22678 18545 22678 4 _0017_
rlabel metal1 s 19412 25126 19412 25126 4 _0018_
rlabel metal1 s 17572 21658 17572 21658 4 _0019_
rlabel metal1 s 10534 28084 10534 28084 4 _0020_
rlabel metal1 s 15962 3400 15962 3400 4 _0021_
rlabel metal1 s 12788 3162 12788 3162 4 _0022_
rlabel metal1 s 9430 3094 9430 3094 4 _0023_
rlabel metal1 s 9062 12410 9062 12410 4 _0024_
rlabel metal1 s 15272 3638 15272 3638 4 _0025_
rlabel metal1 s 10626 3400 10626 3400 4 _0026_
rlabel metal1 s 13248 20502 13248 20502 4 _0027_
rlabel metal1 s 9292 24378 9292 24378 4 _0028_
rlabel metal1 s 11362 30770 11362 30770 4 _0029_
rlabel metal1 s 18262 30260 18262 30260 4 _0030_
rlabel metal1 s 18538 31382 18538 31382 4 _0031_
rlabel metal1 s 18998 30838 18998 30838 4 _0032_
rlabel metal1 s 15732 30362 15732 30362 4 _0033_
rlabel metal1 s 16744 21930 16744 21930 4 _0034_
rlabel metal1 s 16652 22542 16652 22542 4 _0035_
rlabel metal1 s 17572 24378 17572 24378 4 _0036_
rlabel metal1 s 16422 23018 16422 23018 4 _0037_
rlabel metal1 s 14750 14314 14750 14314 4 _0038_
rlabel metal1 s 14439 9622 14439 9622 4 _0039_
rlabel metal1 s 11576 9622 11576 9622 4 _0040_
rlabel metal1 s 10483 10710 10483 10710 4 _0041_
rlabel metal1 s 13830 17238 13830 17238 4 _0042_
rlabel metal2 s 10069 16558 10069 16558 4 _0043_
rlabel metal1 s 11270 24922 11270 24922 4 _0044_
rlabel metal2 s 10442 21726 10442 21726 4 _0045_
rlabel metal2 s 26169 13226 26169 13226 4 _0046_
rlabel metal1 s 26772 10778 26772 10778 4 _0047_
rlabel metal1 s 22080 12614 22080 12614 4 _0048_
rlabel metal1 s 19136 11322 19136 11322 4 _0049_
rlabel metal2 s 22494 18853 22494 18853 4 _0050_
rlabel metal1 s 28208 14994 28208 14994 4 _0051_
rlabel metal1 s 26128 25126 26128 25126 4 _0052_
rlabel metal2 s 26353 19822 26353 19822 4 _0053_
rlabel metal1 s 28826 12886 28826 12886 4 _0054_
rlabel metal1 s 29660 8942 29660 8942 4 _0055_
rlabel metal1 s 24472 10166 24472 10166 4 _0056_
rlabel metal1 s 19913 8874 19913 8874 4 _0057_
rlabel metal1 s 26940 18666 26940 18666 4 _0058_
rlabel metal1 s 30033 16558 30033 16558 4 _0059_
rlabel metal2 s 30318 23698 30318 23698 4 _0060_
rlabel metal1 s 30743 20502 30743 20502 4 _0061_
rlabel metal1 s 12634 13226 12634 13226 4 _0062_
rlabel metal2 s 14030 6562 14030 6562 4 _0063_
rlabel metal2 s 10718 7378 10718 7378 4 _0064_
rlabel metal1 s 9236 7378 9236 7378 4 _0065_
rlabel metal2 s 14306 18054 14306 18054 4 _0066_
rlabel metal1 s 9000 15402 9000 15402 4 _0067_
rlabel metal1 s 9292 27098 9292 27098 4 _0068_
rlabel metal1 s 8464 21862 8464 21862 4 _0069_
rlabel metal1 s 16238 11254 16238 11254 4 _0070_
rlabel metal1 s 14296 11118 14296 11118 4 _0071_
rlabel metal1 s 7406 9146 7406 9146 4 _0072_
rlabel metal1 s 8091 11050 8091 11050 4 _0073_
rlabel metal1 s 14842 18666 14842 18666 4 _0074_
rlabel metal2 s 7309 17646 7309 17646 4 _0075_
rlabel metal2 s 7774 25058 7774 25058 4 _0076_
rlabel metal2 s 7314 22406 7314 22406 4 _0077_
rlabel metal1 s 18988 14994 18988 14994 4 _0078_
rlabel metal1 s 26158 7786 26158 7786 4 _0079_
rlabel metal1 s 21873 7514 21873 7514 4 _0080_
rlabel metal2 s 16877 7854 16877 7854 4 _0081_
rlabel metal2 s 18262 16966 18262 16966 4 _0082_
rlabel metal1 s 25499 16150 25499 16150 4 _0083_
rlabel metal1 s 28566 27064 28566 27064 4 _0084_
rlabel metal2 s 26261 23018 26261 23018 4 _0085_
rlabel metal1 s 28090 13226 28090 13226 4 _0086_
rlabel metal1 s 29164 9146 29164 9146 4 _0087_
rlabel metal1 s 23588 9554 23588 9554 4 _0088_
rlabel metal1 s 18982 9622 18982 9622 4 _0089_
rlabel metal2 s 25801 18666 25801 18666 4 _0090_
rlabel metal1 s 30605 17238 30605 17238 4 _0091_
rlabel metal1 s 29516 24106 29516 24106 4 _0092_
rlabel metal2 s 30686 20910 30686 20910 4 _0093_
rlabel metal2 s 13574 13974 13574 13974 4 _0094_
rlabel metal1 s 13156 4794 13156 4794 4 _0095_
rlabel metal1 s 7401 4182 7401 4182 4 _0096_
rlabel metal1 s 8689 4522 8689 4522 4 _0097_
rlabel metal1 s 11955 19414 11955 19414 4 _0098_
rlabel metal2 s 7038 14178 7038 14178 4 _0099_
rlabel metal1 s 7222 26010 7222 26010 4 _0100_
rlabel metal2 s 7309 19822 7309 19822 4 _0101_
rlabel metal1 s 24456 13226 24456 13226 4 _0102_
rlabel metal1 s 25571 11050 25571 11050 4 _0103_
rlabel metal1 s 21558 12138 21558 12138 4 _0104_
rlabel metal1 s 18032 11322 18032 11322 4 _0105_
rlabel metal1 s 20787 19414 20787 19414 4 _0106_
rlabel metal2 s 26537 15402 26537 15402 4 _0107_
rlabel metal1 s 23966 26214 23966 26214 4 _0108_
rlabel metal1 s 24012 20026 24012 20026 4 _0109_
rlabel metal2 s 21394 14382 21394 14382 4 _0110_
rlabel metal1 s 24364 5610 24364 5610 4 _0111_
rlabel metal1 s 21201 4590 21201 4590 4 _0112_
rlabel metal1 s 17848 4794 17848 4794 4 _0113_
rlabel metal1 s 19442 18666 19442 18666 4 _0114_
rlabel metal1 s 21666 16184 21666 16184 4 _0115_
rlabel metal1 s 23368 26214 23368 26214 4 _0116_
rlabel metal2 s 23506 21794 23506 21794 4 _0117_
rlabel metal1 s 10902 14042 10902 14042 4 _0118_
rlabel metal2 s 11725 5610 11725 5610 4 _0119_
rlabel metal2 s 5934 6562 5934 6562 4 _0120_
rlabel metal1 s 6424 6358 6424 6358 4 _0121_
rlabel metal2 s 10626 19142 10626 19142 4 _0122_
rlabel metal2 s 6026 14178 6026 14178 4 _0123_
rlabel metal2 s 7590 26112 7590 26112 4 _0124_
rlabel metal1 s 6568 19346 6568 19346 4 _0125_
rlabel metal1 s 2663 13974 2663 13974 4 _0126_
rlabel metal1 s 6757 11798 6757 11798 4 _0127_
rlabel metal1 s 2852 9146 2852 9146 4 _0128_
rlabel metal1 s 2336 11118 2336 11118 4 _0129_
rlabel metal1 s 3542 18870 3542 18870 4 _0130_
rlabel metal1 s 3848 16490 3848 16490 4 _0131_
rlabel metal1 s 4411 24854 4411 24854 4 _0132_
rlabel metal1 s 4048 22950 4048 22950 4 _0133_
rlabel metal2 s 18625 13974 18625 13974 4 _0134_
rlabel metal1 s 23874 5882 23874 5882 4 _0135_
rlabel metal1 s 20086 5270 20086 5270 4 _0136_
rlabel metal1 s 17250 5338 17250 5338 4 _0137_
rlabel metal2 s 17521 19414 17521 19414 4 _0138_
rlabel metal2 s 22121 16558 22121 16558 4 _0139_
rlabel metal2 s 23133 27438 23133 27438 4 _0140_
rlabel metal1 s 23455 22678 23455 22678 4 _0141_
rlabel metal1 s 3542 13498 3542 13498 4 _0142_
rlabel metal1 s 6869 11050 6869 11050 4 _0143_
rlabel metal2 s 2622 10438 2622 10438 4 _0144_
rlabel metal1 s 3675 11730 3675 11730 4 _0145_
rlabel metal2 s 3082 19142 3082 19142 4 _0146_
rlabel metal1 s 3450 16762 3450 16762 4 _0147_
rlabel metal1 s 5106 24922 5106 24922 4 _0148_
rlabel metal1 s 3710 22678 3710 22678 4 _0149_
rlabel metal2 s 17613 14994 17613 14994 4 _0150_
rlabel metal1 s 28704 7514 28704 7514 4 _0151_
rlabel metal1 s 20000 7378 20000 7378 4 _0152_
rlabel metal1 s 16872 8466 16872 8466 4 _0153_
rlabel metal1 s 17418 18326 17418 18326 4 _0154_
rlabel metal1 s 24364 16490 24364 16490 4 _0155_
rlabel metal2 s 26353 27438 26353 27438 4 _0156_
rlabel metal1 s 27917 23018 27917 23018 4 _0157_
rlabel metal2 s 12466 14824 12466 14824 4 _0158_
rlabel metal2 s 13468 7378 13468 7378 4 _0159_
rlabel metal2 s 5658 7650 5658 7650 4 _0160_
rlabel metal1 s 5791 6698 5791 6698 4 _0161_
rlabel metal2 s 11914 18530 11914 18530 4 _0162_
rlabel metal1 s 6992 16762 6992 16762 4 _0163_
rlabel metal1 s 8954 28458 8954 28458 4 _0164_
rlabel metal2 s 6210 21318 6210 21318 4 _0165_
rlabel metal1 s 20286 27574 20286 27574 4 _0166_
rlabel metal1 s 20700 27302 20700 27302 4 _0167_
rlabel metal1 s 20884 27438 20884 27438 4 _0168_
rlabel metal1 s 21022 27098 21022 27098 4 _0169_
rlabel metal1 s 14490 26894 14490 26894 4 _0170_
rlabel metal1 s 14076 26962 14076 26962 4 _0171_
rlabel metal1 s 10580 24242 10580 24242 4 _0172_
rlabel metal1 s 22494 23086 22494 23086 4 _0173_
rlabel metal2 s 20102 24582 20102 24582 4 _0174_
rlabel metal2 s 12558 16524 12558 16524 4 _0175_
rlabel metal2 s 20378 24004 20378 24004 4 _0176_
rlabel metal2 s 15318 23868 15318 23868 4 _0177_
rlabel metal1 s 15134 23494 15134 23494 4 _0178_
rlabel metal1 s 20562 23086 20562 23086 4 _0179_
rlabel metal1 s 20884 22406 20884 22406 4 _0180_
rlabel metal1 s 15134 23732 15134 23732 4 _0181_
rlabel metal2 s 15502 23290 15502 23290 4 _0182_
rlabel metal1 s 19642 23154 19642 23154 4 _0183_
rlabel metal1 s 16146 23834 16146 23834 4 _0184_
rlabel metal1 s 14490 22746 14490 22746 4 _0185_
rlabel metal2 s 16146 22039 16146 22039 4 _0186_
rlabel metal1 s 16100 22066 16100 22066 4 _0187_
rlabel metal1 s 13984 29614 13984 29614 4 _0188_
rlabel metal1 s 13938 29138 13938 29138 4 _0189_
rlabel metal1 s 16744 26962 16744 26962 4 _0190_
rlabel metal1 s 14582 28050 14582 28050 4 _0191_
rlabel metal1 s 15594 29818 15594 29818 4 _0192_
rlabel metal1 s 13800 30294 13800 30294 4 _0193_
rlabel metal1 s 16238 30158 16238 30158 4 _0194_
rlabel metal1 s 18354 30736 18354 30736 4 _0195_
rlabel metal1 s 17894 30192 17894 30192 4 _0196_
rlabel metal1 s 18032 31314 18032 31314 4 _0197_
rlabel metal1 s 24426 22440 24426 22440 4 _0198_
rlabel metal2 s 21298 9826 21298 9826 4 _0199_
rlabel metal1 s 21735 21862 21735 21862 4 _0200_
rlabel metal1 s 28290 20026 28290 20026 4 _0201_
rlabel metal1 s 22954 24140 22954 24140 4 _0202_
rlabel metal1 s 23230 23732 23230 23732 4 _0203_
rlabel metal1 s 26818 21114 26818 21114 4 _0204_
rlabel metal1 s 26910 22610 26910 22610 4 _0205_
rlabel metal1 s 25346 22576 25346 22576 4 _0206_
rlabel metal1 s 26956 21454 26956 21454 4 _0207_
rlabel metal1 s 24472 24650 24472 24650 4 _0208_
rlabel metal1 s 24288 24718 24288 24718 4 _0209_
rlabel metal1 s 25852 21522 25852 21522 4 _0210_
rlabel metal2 s 17342 21590 17342 21590 4 _0211_
rlabel metal1 s 8050 24106 8050 24106 4 _0212_
rlabel metal1 s 6394 23018 6394 23018 4 _0213_
rlabel metal1 s 5980 23018 5980 23018 4 _0214_
rlabel metal1 s 7176 22950 7176 22950 4 _0215_
rlabel metal1 s 8188 21930 8188 21930 4 _0216_
rlabel metal2 s 10168 25874 10168 25874 4 _0217_
rlabel metal1 s 14030 24106 14030 24106 4 _0218_
rlabel metal1 s 10304 25398 10304 25398 4 _0219_
rlabel metal2 s 10074 24480 10074 24480 4 _0220_
rlabel metal1 s 9108 20298 9108 20298 4 _0221_
rlabel metal1 s 9890 22134 9890 22134 4 _0222_
rlabel metal2 s 12190 23256 12190 23256 4 _0223_
rlabel metal1 s 9890 22032 9890 22032 4 _0224_
rlabel metal1 s 10258 22202 10258 22202 4 _0225_
rlabel metal1 s 9614 24174 9614 24174 4 _0226_
rlabel metal2 s 26082 24004 26082 24004 4 _0227_
rlabel metal2 s 25990 24480 25990 24480 4 _0228_
rlabel metal1 s 27002 24310 27002 24310 4 _0229_
rlabel metal1 s 25300 24174 25300 24174 4 _0230_
rlabel metal1 s 11983 24174 11983 24174 4 _0231_
rlabel metal1 s 6509 24310 6509 24310 4 _0232_
rlabel metal1 s 9982 24310 9982 24310 4 _0233_
rlabel metal2 s 9706 25670 9706 25670 4 _0234_
rlabel metal1 s 11408 24174 11408 24174 4 _0235_
rlabel metal1 s 11270 24208 11270 24208 4 _0236_
rlabel metal1 s 12236 24038 12236 24038 4 _0237_
rlabel metal1 s 13478 21590 13478 21590 4 _0238_
rlabel metal1 s 25714 16048 25714 16048 4 _0239_
rlabel metal2 s 26266 15504 26266 15504 4 _0240_
rlabel metal2 s 25806 16524 25806 16524 4 _0241_
rlabel metal1 s 25990 16184 25990 16184 4 _0242_
rlabel metal1 s 21574 16150 21574 16150 4 _0243_
rlabel metal1 s 9062 17238 9062 17238 4 _0244_
rlabel metal1 s 9936 16014 9936 16014 4 _0245_
rlabel metal1 s 8648 15674 8648 15674 4 _0246_
rlabel metal1 s 9844 15946 9844 15946 4 _0247_
rlabel metal1 s 9982 16116 9982 16116 4 _0248_
rlabel metal1 s 10534 15878 10534 15878 4 _0249_
rlabel metal1 s 10074 3604 10074 3604 4 _0250_
rlabel metal2 s 24886 18870 24886 18870 4 _0251_
rlabel metal1 s 21482 18122 21482 18122 4 _0252_
rlabel metal1 s 20562 17782 20562 17782 4 _0253_
rlabel metal1 s 21114 17850 21114 17850 4 _0254_
rlabel metal1 s 16238 17680 16238 17680 4 _0255_
rlabel metal1 s 15134 19278 15134 19278 4 _0256_
rlabel metal1 s 15824 17782 15824 17782 4 _0257_
rlabel metal1 s 13018 17850 13018 17850 4 _0258_
rlabel metal1 s 16422 17816 16422 17816 4 _0259_
rlabel metal1 s 16422 17306 16422 17306 4 _0260_
rlabel metal1 s 15778 17714 15778 17714 4 _0261_
rlabel metal1 s 15134 3604 15134 3604 4 _0262_
rlabel metal1 s 20608 10234 20608 10234 4 _0263_
rlabel metal1 s 19918 10472 19918 10472 4 _0264_
rlabel metal1 s 19412 9146 19412 9146 4 _0265_
rlabel metal2 s 19550 8534 19550 8534 4 _0266_
rlabel metal2 s 20102 10336 20102 10336 4 _0267_
rlabel metal1 s 8602 10642 8602 10642 4 _0268_
rlabel metal1 s 9568 10166 9568 10166 4 _0269_
rlabel metal1 s 9200 6426 9200 6426 4 _0270_
rlabel metal2 s 9890 9282 9890 9282 4 _0271_
rlabel metal1 s 10626 10030 10626 10030 4 _0272_
rlabel metal1 s 10028 10234 10028 10234 4 _0273_
rlabel metal1 s 9384 12206 9384 12206 4 _0274_
rlabel metal1 s 23230 8942 23230 8942 4 _0275_
rlabel metal2 s 22862 10234 22862 10234 4 _0276_
rlabel metal1 s 22632 8602 22632 8602 4 _0277_
rlabel metal1 s 22540 6426 22540 6426 4 _0278_
rlabel metal1 s 17250 8908 17250 8908 4 _0279_
rlabel metal1 s 7084 10642 7084 10642 4 _0280_
rlabel metal1 s 9982 9010 9982 9010 4 _0281_
rlabel metal1 s 8878 7854 8878 7854 4 _0282_
rlabel metal1 s 10534 7718 10534 7718 4 _0283_
rlabel metal1 s 11454 8942 11454 8942 4 _0284_
rlabel metal1 s 10350 4114 10350 4114 4 _0285_
rlabel metal1 s 9706 3604 9706 3604 4 _0286_
rlabel metal1 s 26726 8908 26726 8908 4 _0287_
rlabel metal2 s 26450 10336 26450 10336 4 _0288_
rlabel metal1 s 26450 8602 26450 8602 4 _0289_
rlabel metal1 s 26496 6630 26496 6630 4 _0290_
rlabel metal3 s 14858 8483 14858 8483 4 _0291_
rlabel metal1 s 14398 10064 14398 10064 4 _0292_
rlabel metal2 s 14950 9214 14950 9214 4 _0293_
rlabel metal2 s 13754 7684 13754 7684 4 _0294_
rlabel metal1 s 14812 8398 14812 8398 4 _0295_
rlabel metal1 s 15456 8466 15456 8466 4 _0296_
rlabel metal2 s 14582 6018 14582 6018 4 _0297_
rlabel metal1 s 13294 3060 13294 3060 4 _0298_
rlabel metal1 s 29440 13158 29440 13158 4 _0299_
rlabel metal1 s 23414 13770 23414 13770 4 _0300_
rlabel metal1 s 22034 13940 22034 13940 4 _0301_
rlabel metal1 s 21804 13906 21804 13906 4 _0302_
rlabel metal2 s 22126 13736 22126 13736 4 _0303_
rlabel metal2 s 16606 13566 16606 13566 4 _0304_
rlabel metal1 s 15962 13260 15962 13260 4 _0305_
rlabel metal1 s 13524 12818 13524 12818 4 _0306_
rlabel metal1 s 15134 12954 15134 12954 4 _0307_
rlabel metal2 s 16146 13345 16146 13345 4 _0308_
rlabel metal1 s 15824 4046 15824 4046 4 _0309_
rlabel metal1 s 15410 3570 15410 3570 4 _0310_
rlabel metal2 s 13938 30022 13938 30022 4 _0311_
rlabel metal1 s 14076 29818 14076 29818 4 _0312_
rlabel metal1 s 19366 29648 19366 29648 4 _0313_
rlabel metal1 s 10994 24752 10994 24752 4 _0314_
rlabel metal1 s 21298 13906 21298 13906 4 _0315_
rlabel metal1 s 14720 28186 14720 28186 4 _0316_
rlabel metal1 s 18584 27098 18584 27098 4 _0317_
rlabel metal1 s 14686 26282 14686 26282 4 _0318_
rlabel metal1 s 15180 25942 15180 25942 4 _0319_
rlabel metal1 s 14996 17714 14996 17714 4 _0320_
rlabel metal1 s 14858 14042 14858 14042 4 _0321_
rlabel metal1 s 16008 5542 16008 5542 4 _0322_
rlabel metal1 s 14996 9146 14996 9146 4 _0323_
rlabel metal2 s 12466 8636 12466 8636 4 _0324_
rlabel metal1 s 11546 9146 11546 9146 4 _0325_
rlabel metal1 s 19642 9894 19642 9894 4 _0326_
rlabel metal2 s 11546 10948 11546 10948 4 _0327_
rlabel metal2 s 21666 19244 21666 19244 4 _0328_
rlabel metal1 s 13570 17170 13570 17170 4 _0329_
rlabel metal1 s 15548 15878 15548 15878 4 _0330_
rlabel metal1 s 10580 16218 10580 16218 4 _0331_
rlabel metal1 s 24426 25126 24426 25126 4 _0332_
rlabel metal1 s 11454 24786 11454 24786 4 _0333_
rlabel metal1 s 8970 22610 8970 22610 4 _0334_
rlabel metal2 s 10626 21556 10626 21556 4 _0335_
rlabel metal2 s 18170 26571 18170 26571 4 _0336_
rlabel metal2 s 25622 25874 25622 25874 4 _0337_
rlabel metal1 s 26680 12954 26680 12954 4 _0338_
rlabel metal1 s 26772 10642 26772 10642 4 _0339_
rlabel metal1 s 22586 12818 22586 12818 4 _0340_
rlabel metal1 s 18952 11118 18952 11118 4 _0341_
rlabel metal1 s 21206 18734 21206 18734 4 _0342_
rlabel metal1 s 28658 15504 28658 15504 4 _0343_
rlabel metal1 s 26082 25364 26082 25364 4 _0344_
rlabel metal1 s 26772 20434 26772 20434 4 _0345_
rlabel metal1 s 16158 27030 16158 27030 4 _0346_
rlabel metal1 s 19458 25942 19458 25942 4 _0347_
rlabel metal1 s 25438 25772 25438 25772 4 _0348_
rlabel metal1 s 29026 12614 29026 12614 4 _0349_
rlabel metal1 s 29348 10030 29348 10030 4 _0350_
rlabel metal1 s 24058 10030 24058 10030 4 _0351_
rlabel metal2 s 20378 10166 20378 10166 4 _0352_
rlabel metal1 s 26726 18054 26726 18054 4 _0353_
rlabel metal1 s 30590 17646 30590 17646 4 _0354_
rlabel metal2 s 29394 24582 29394 24582 4 _0355_
rlabel metal1 s 31234 21012 31234 21012 4 _0356_
rlabel metal1 s 13984 27438 13984 27438 4 _0357_
rlabel metal2 s 9752 23868 9752 23868 4 _0358_
rlabel metal1 s 13271 13498 13271 13498 4 _0359_
rlabel metal1 s 14260 6290 14260 6290 4 _0360_
rlabel metal1 s 10534 6732 10534 6732 4 _0361_
rlabel metal1 s 9154 6970 9154 6970 4 _0362_
rlabel metal1 s 14030 17646 14030 17646 4 _0363_
rlabel metal1 s 8740 15130 8740 15130 4 _0364_
rlabel metal1 s 9476 26962 9476 26962 4 _0365_
rlabel metal2 s 8970 21556 8970 21556 4 _0366_
rlabel metal1 s 15054 27030 15054 27030 4 _0367_
rlabel metal2 s 15410 26350 15410 26350 4 _0368_
rlabel metal1 s 9154 22542 9154 22542 4 _0369_
rlabel metal1 s 16514 11152 16514 11152 4 _0370_
rlabel metal2 s 14214 11254 14214 11254 4 _0371_
rlabel metal1 s 7820 8942 7820 8942 4 _0372_
rlabel metal1 s 8832 10778 8832 10778 4 _0373_
rlabel metal1 s 14812 18394 14812 18394 4 _0374_
rlabel metal1 s 7774 18258 7774 18258 4 _0375_
rlabel metal1 s 8004 24786 8004 24786 4 _0376_
rlabel metal2 s 8050 22304 8050 22304 4 _0377_
rlabel metal1 s 17664 27098 17664 27098 4 _0378_
rlabel metal1 s 25070 26316 25070 26316 4 _0379_
rlabel metal1 s 18722 14586 18722 14586 4 _0380_
rlabel metal1 s 26404 7514 26404 7514 4 _0381_
rlabel metal1 s 21574 7378 21574 7378 4 _0382_
rlabel metal1 s 16468 8466 16468 8466 4 _0383_
rlabel metal1 s 18722 16558 18722 16558 4 _0384_
rlabel metal1 s 25898 16558 25898 16558 4 _0385_
rlabel metal1 s 28382 26554 28382 26554 4 _0386_
rlabel metal1 s 26864 21862 26864 21862 4 _0387_
rlabel metal1 s 18584 25874 18584 25874 4 _0388_
rlabel metal1 s 25438 25296 25438 25296 4 _0389_
rlabel metal1 s 27830 13294 27830 13294 4 _0390_
rlabel metal1 s 28888 8942 28888 8942 4 _0391_
rlabel metal1 s 23782 9146 23782 9146 4 _0392_
rlabel metal1 s 18630 9452 18630 9452 4 _0393_
rlabel metal2 s 25990 18870 25990 18870 4 _0394_
rlabel metal1 s 31004 17170 31004 17170 4 _0395_
rlabel metal1 s 28382 24242 28382 24242 4 _0396_
rlabel metal1 s 30452 21522 30452 21522 4 _0397_
rlabel metal1 s 14030 26010 14030 26010 4 _0398_
rlabel metal2 s 14490 13821 14490 13821 4 _0399_
rlabel metal1 s 13846 14042 13846 14042 4 _0400_
rlabel metal1 s 13386 4624 13386 4624 4 _0401_
rlabel metal1 s 7222 4590 7222 4590 4 _0402_
rlabel metal1 s 9890 4624 9890 4624 4 _0403_
rlabel metal1 s 12236 18394 12236 18394 4 _0404_
rlabel metal1 s 7406 13906 7406 13906 4 _0405_
rlabel metal1 s 7498 25908 7498 25908 4 _0406_
rlabel metal1 s 7682 19482 7682 19482 4 _0407_
rlabel metal1 s 14741 27540 14741 27540 4 _0408_
rlabel metal1 s 19044 26350 19044 26350 4 _0409_
rlabel metal1 s 25116 25330 25116 25330 4 _0410_
rlabel metal1 s 24288 12954 24288 12954 4 _0411_
rlabel metal1 s 25760 10778 25760 10778 4 _0412_
rlabel metal1 s 21620 11322 21620 11322 4 _0413_
rlabel metal1 s 18262 11152 18262 11152 4 _0414_
rlabel metal2 s 21206 19380 21206 19380 4 _0415_
rlabel metal2 s 26174 15878 26174 15878 4 _0416_
rlabel metal1 s 24058 25466 24058 25466 4 _0417_
rlabel metal1 s 24702 19822 24702 19822 4 _0418_
rlabel metal1 s 19274 26282 19274 26282 4 _0419_
rlabel metal1 s 23076 25330 23076 25330 4 _0420_
rlabel metal1 s 21482 13804 21482 13804 4 _0421_
rlabel metal1 s 24656 6426 24656 6426 4 _0422_
rlabel metal1 s 21436 5202 21436 5202 4 _0423_
rlabel metal1 s 18216 4590 18216 4590 4 _0424_
rlabel metal1 s 19090 19346 19090 19346 4 _0425_
rlabel metal1 s 21482 15980 21482 15980 4 _0426_
rlabel metal2 s 23506 25908 23506 25908 4 _0427_
rlabel metal1 s 24426 21896 24426 21896 4 _0428_
rlabel metal1 s 13386 26384 13386 26384 4 _0429_
rlabel metal1 s 6578 25772 6578 25772 4 _0430_
rlabel metal1 s 11362 13906 11362 13906 4 _0431_
rlabel metal1 s 11960 6290 11960 6290 4 _0432_
rlabel metal1 s 5980 5882 5980 5882 4 _0433_
rlabel metal1 s 6624 6290 6624 6290 4 _0434_
rlabel metal1 s 10856 18734 10856 18734 4 _0435_
rlabel metal1 s 6302 13906 6302 13906 4 _0436_
rlabel metal1 s 7774 25840 7774 25840 4 _0437_
rlabel metal1 s 6348 18938 6348 18938 4 _0438_
rlabel metal1 s 9752 27030 9752 27030 4 _0439_
rlabel metal1 s 5888 22134 5888 22134 4 _0440_
rlabel metal1 s 2990 14994 2990 14994 4 _0441_
rlabel metal1 s 7176 10778 7176 10778 4 _0442_
rlabel metal1 s 3450 8942 3450 8942 4 _0443_
rlabel metal1 s 1978 11084 1978 11084 4 _0444_
rlabel metal1 s 2990 18734 2990 18734 4 _0445_
rlabel metal1 s 3864 16218 3864 16218 4 _0446_
rlabel metal2 s 5474 25602 5474 25602 4 _0447_
rlabel metal1 s 5014 22202 5014 22202 4 _0448_
rlabel metal1 s 18170 26350 18170 26350 4 _0449_
rlabel metal1 s 24610 26894 24610 26894 4 _0450_
rlabel metal1 s 17802 14280 17802 14280 4 _0451_
rlabel metal1 s 24196 5678 24196 5678 4 _0452_
rlabel metal1 s 19734 5202 19734 5202 4 _0453_
rlabel metal1 s 17388 5202 17388 5202 4 _0454_
rlabel metal1 s 17664 18938 17664 18938 4 _0455_
rlabel metal1 s 22586 15674 22586 15674 4 _0456_
rlabel metal1 s 23368 27098 23368 27098 4 _0457_
rlabel metal1 s 24150 22746 24150 22746 4 _0458_
rlabel metal2 s 9154 26962 9154 26962 4 _0459_
rlabel metal1 s 5658 22576 5658 22576 4 _0460_
rlabel metal1 s 3910 13294 3910 13294 4 _0461_
rlabel metal1 s 7176 11118 7176 11118 4 _0462_
rlabel metal1 s 3404 10030 3404 10030 4 _0463_
rlabel metal1 s 4784 11866 4784 11866 4 _0464_
rlabel metal1 s 3542 18734 3542 18734 4 _0465_
rlabel metal1 s 3174 16524 3174 16524 4 _0466_
rlabel metal1 s 5566 24854 5566 24854 4 _0467_
rlabel metal1 s 3358 22508 3358 22508 4 _0468_
rlabel metal1 s 18584 26962 18584 26962 4 _0469_
rlabel metal2 s 27922 22916 27922 22916 4 _0470_
rlabel metal1 s 17848 14586 17848 14586 4 _0471_
rlabel metal1 s 28198 7378 28198 7378 4 _0472_
rlabel metal1 s 19596 7378 19596 7378 4 _0473_
rlabel metal1 s 16054 8500 16054 8500 4 _0474_
rlabel metal1 s 17066 18224 17066 18224 4 _0475_
rlabel metal1 s 24058 16762 24058 16762 4 _0476_
rlabel metal1 s 26818 27098 26818 27098 4 _0477_
rlabel metal1 s 28290 22746 28290 22746 4 _0478_
rlabel metal1 s 13386 28084 13386 28084 4 _0479_
rlabel metal1 s 9338 27948 9338 27948 4 _0480_
rlabel metal1 s 12696 14382 12696 14382 4 _0481_
rlabel metal1 s 13570 7786 13570 7786 4 _0482_
rlabel metal1 s 6302 7378 6302 7378 4 _0483_
rlabel metal1 s 6210 7514 6210 7514 4 _0484_
rlabel metal2 s 13018 18700 13018 18700 4 _0485_
rlabel metal1 s 7176 16558 7176 16558 4 _0486_
rlabel metal1 s 8648 28186 8648 28186 4 _0487_
rlabel metal1 s 6394 21012 6394 21012 4 _0488_
rlabel metal3 s 28336 31892 28336 31892 4 clk
rlabel metal2 s 20516 12716 20516 12716 4 clknet_0_clk
rlabel metal1 s 10350 3468 10350 3468 4 clknet_4_0_0_clk
rlabel metal1 s 25990 11118 25990 11118 4 clknet_4_10_0_clk
rlabel metal1 s 28520 14994 28520 14994 4 clknet_4_11_0_clk
rlabel metal1 s 20148 19346 20148 19346 4 clknet_4_12_0_clk
rlabel metal1 s 23138 22644 23138 22644 4 clknet_4_13_0_clk
rlabel metal1 s 30636 20434 30636 20434 4 clknet_4_14_0_clk
rlabel metal1 s 30590 23732 30590 23732 4 clknet_4_15_0_clk
rlabel metal1 s 2300 14382 2300 14382 4 clknet_4_1_0_clk
rlabel metal1 s 16652 7854 16652 7854 4 clknet_4_2_0_clk
rlabel metal1 s 13984 13838 13984 13838 4 clknet_4_3_0_clk
rlabel metal1 s 2530 19380 2530 19380 4 clknet_4_4_0_clk
rlabel metal2 s 4002 25772 4002 25772 4 clknet_4_5_0_clk
rlabel metal1 s 14582 18122 14582 18122 4 clknet_4_6_0_clk
rlabel metal1 s 10810 31212 10810 31212 4 clknet_4_7_0_clk
rlabel metal1 s 19918 5236 19918 5236 4 clknet_4_8_0_clk
rlabel metal1 s 21436 12750 21436 12750 4 clknet_4_9_0_clk
rlabel metal3 s 820 30668 820 30668 4 data_in[0]
rlabel metal2 s 29026 823 29026 823 4 data_in[1]
rlabel metal3 s 820 6188 820 6188 4 data_in[2]
rlabel metal3 s 820 18428 820 18428 4 data_in[3]
rlabel metal1 s 7176 32402 7176 32402 4 data_in[4]
rlabel metal1 s 12972 32402 12972 32402 4 data_in[5]
rlabel metal1 s 30360 32402 30360 32402 4 data_in[6]
rlabel metal1 s 31648 7786 31648 7786 4 data_in[7]
rlabel metal2 s 23230 1095 23230 1095 4 data_out[0]
rlabel metal2 s 46 1554 46 1554 4 data_out[1]
rlabel metal2 s 5842 1520 5842 1520 4 data_out[2]
rlabel metal3 s 1096 12308 1096 12308 4 data_out[3]
rlabel metal2 s 31418 1853 31418 1853 4 data_out[4]
rlabel metal2 s 11638 1520 11638 1520 4 data_out[5]
rlabel metal1 s 31648 20026 31648 20026 4 data_out[6]
rlabel metal3 s 31886 25908 31886 25908 4 data_out[7]
rlabel metal1 s 19090 32538 19090 32538 4 empty
rlabel metal1 s 24748 32538 24748 32538 4 error
rlabel metal1 s 16376 14518 16376 14518 4 fifo\[0\]\[0\]
rlabel metal1 s 15640 9486 15640 9486 4 fifo\[0\]\[1\]
rlabel metal2 s 12926 9860 12926 9860 4 fifo\[0\]\[2\]
rlabel metal2 s 11362 10982 11362 10982 4 fifo\[0\]\[3\]
rlabel metal1 s 16146 17272 16146 17272 4 fifo\[0\]\[4\]
rlabel metal1 s 11822 16660 11822 16660 4 fifo\[0\]\[5\]
rlabel metal1 s 12190 25364 12190 25364 4 fifo\[0\]\[6\]
rlabel metal1 s 11086 21658 11086 21658 4 fifo\[0\]\[7\]
rlabel metal2 s 12834 13532 12834 13532 4 fifo\[10\]\[0\]
rlabel metal1 s 13110 6222 13110 6222 4 fifo\[10\]\[1\]
rlabel metal2 s 8326 7480 8326 7480 4 fifo\[10\]\[2\]
rlabel metal2 s 8602 6800 8602 6800 4 fifo\[10\]\[3\]
rlabel metal1 s 11546 19482 11546 19482 4 fifo\[10\]\[4\]
rlabel metal2 s 7222 15028 7222 15028 4 fifo\[10\]\[5\]
rlabel metal1 s 10258 25296 10258 25296 4 fifo\[10\]\[6\]
rlabel metal2 s 7774 19822 7774 19822 4 fifo\[10\]\[7\]
rlabel metal1 s 4370 13974 4370 13974 4 fifo\[11\]\[0\]
rlabel metal1 s 8142 11832 8142 11832 4 fifo\[11\]\[1\]
rlabel metal1 s 4968 10030 4968 10030 4 fifo\[11\]\[2\]
rlabel metal1 s 4968 11118 4968 11118 4 fifo\[11\]\[3\]
rlabel metal1 s 5474 19482 5474 19482 4 fifo\[11\]\[4\]
rlabel metal1 s 6026 16626 6026 16626 4 fifo\[11\]\[5\]
rlabel metal2 s 6946 24956 6946 24956 4 fifo\[11\]\[6\]
rlabel metal1 s 6210 20978 6210 20978 4 fifo\[11\]\[7\]
rlabel metal2 s 19734 14722 19734 14722 4 fifo\[12\]\[0\]
rlabel metal1 s 25668 6766 25668 6766 4 fifo\[12\]\[1\]
rlabel metal2 s 21574 5644 21574 5644 4 fifo\[12\]\[2\]
rlabel metal1 s 18446 6222 18446 6222 4 fifo\[12\]\[3\]
rlabel metal1 s 19734 19890 19734 19890 4 fifo\[12\]\[4\]
rlabel metal1 s 23322 16116 23322 16116 4 fifo\[12\]\[5\]
rlabel metal1 s 24610 27438 24610 27438 4 fifo\[12\]\[6\]
rlabel metal1 s 24656 22406 24656 22406 4 fifo\[12\]\[7\]
rlabel metal1 s 4094 13906 4094 13906 4 fifo\[13\]\[0\]
rlabel metal1 s 6072 11662 6072 11662 4 fifo\[13\]\[1\]
rlabel metal1 s 5382 10540 5382 10540 4 fifo\[13\]\[2\]
rlabel metal1 s 4462 12206 4462 12206 4 fifo\[13\]\[3\]
rlabel metal2 s 5198 19142 5198 19142 4 fifo\[13\]\[4\]
rlabel metal1 s 5244 17646 5244 17646 4 fifo\[13\]\[5\]
rlabel metal1 s 5704 25398 5704 25398 4 fifo\[13\]\[6\]
rlabel metal1 s 5336 23086 5336 23086 4 fifo\[13\]\[7\]
rlabel metal1 s 20010 15470 20010 15470 4 fifo\[14\]\[0\]
rlabel metal1 s 27324 8058 27324 8058 4 fifo\[14\]\[1\]
rlabel metal1 s 21758 7208 21758 7208 4 fifo\[14\]\[2\]
rlabel metal1 s 18354 8908 18354 8908 4 fifo\[14\]\[3\]
rlabel metal1 s 18814 18054 18814 18054 4 fifo\[14\]\[4\]
rlabel metal2 s 25898 16932 25898 16932 4 fifo\[14\]\[5\]
rlabel metal1 s 27370 27302 27370 27302 4 fifo\[14\]\[6\]
rlabel metal1 s 28658 22950 28658 22950 4 fifo\[14\]\[7\]
rlabel metal1 s 13524 14790 13524 14790 4 fifo\[15\]\[0\]
rlabel metal1 s 14352 7514 14352 7514 4 fifo\[15\]\[1\]
rlabel metal1 s 8142 7956 8142 7956 4 fifo\[15\]\[2\]
rlabel metal1 s 7038 8398 7038 8398 4 fifo\[15\]\[3\]
rlabel metal1 s 13800 18938 13800 18938 4 fifo\[15\]\[4\]
rlabel metal1 s 8878 17102 8878 17102 4 fifo\[15\]\[5\]
rlabel metal2 s 9872 25874 9872 25874 4 fifo\[15\]\[6\]
rlabel metal1 s 7222 21930 7222 21930 4 fifo\[15\]\[7\]
rlabel metal2 s 27278 13736 27278 13736 4 fifo\[1\]\[0\]
rlabel metal2 s 28106 11492 28106 11492 4 fifo\[1\]\[1\]
rlabel metal1 s 23552 11866 23552 11866 4 fifo\[1\]\[2\]
rlabel metal1 s 20838 11526 20838 11526 4 fifo\[1\]\[3\]
rlabel metal2 s 23046 18683 23046 18683 4 fifo\[1\]\[4\]
rlabel metal1 s 27462 15130 27462 15130 4 fifo\[1\]\[5\]
rlabel metal1 s 25714 24752 25714 24752 4 fifo\[1\]\[6\]
rlabel metal1 s 27370 20026 27370 20026 4 fifo\[1\]\[7\]
rlabel metal1 s 29946 12954 29946 12954 4 fifo\[2\]\[0\]
rlabel metal1 s 30912 9554 30912 9554 4 fifo\[2\]\[1\]
rlabel metal1 s 26174 9350 26174 9350 4 fifo\[2\]\[2\]
rlabel metal1 s 21298 9010 21298 9010 4 fifo\[2\]\[3\]
rlabel metal1 s 28198 18938 28198 18938 4 fifo\[2\]\[4\]
rlabel metal1 s 30958 16490 30958 16490 4 fifo\[2\]\[5\]
rlabel metal2 s 28750 24208 28750 24208 4 fifo\[2\]\[6\]
rlabel metal1 s 29716 20570 29716 20570 4 fifo\[2\]\[7\]
rlabel metal1 s 14720 13430 14720 13430 4 fifo\[3\]\[0\]
rlabel metal2 s 15502 7752 15502 7752 4 fifo\[3\]\[1\]
rlabel metal2 s 9798 8500 9798 8500 4 fifo\[3\]\[2\]
rlabel metal1 s 10212 7514 10212 7514 4 fifo\[3\]\[3\]
rlabel metal1 s 13570 18054 13570 18054 4 fifo\[3\]\[4\]
rlabel metal1 s 9844 15674 9844 15674 4 fifo\[3\]\[5\]
rlabel metal1 s 10258 27302 10258 27302 4 fifo\[3\]\[6\]
rlabel metal1 s 8740 20434 8740 20434 4 fifo\[3\]\[7\]
rlabel metal1 s 16238 13158 16238 13158 4 fifo\[4\]\[0\]
rlabel metal2 s 15502 10540 15502 10540 4 fifo\[4\]\[1\]
rlabel metal2 s 8418 10234 8418 10234 4 fifo\[4\]\[2\]
rlabel metal1 s 9660 11254 9660 11254 4 fifo\[4\]\[3\]
rlabel metal1 s 16054 18938 16054 18938 4 fifo\[4\]\[4\]
rlabel metal1 s 8832 17850 8832 17850 4 fifo\[4\]\[5\]
rlabel metal1 s 8648 25126 8648 25126 4 fifo\[4\]\[6\]
rlabel metal2 s 7958 22916 7958 22916 4 fifo\[4\]\[7\]
rlabel metal1 s 20194 14892 20194 14892 4 fifo\[5\]\[0\]
rlabel metal1 s 27416 7718 27416 7718 4 fifo\[5\]\[1\]
rlabel metal1 s 22011 8466 22011 8466 4 fifo\[5\]\[2\]
rlabel metal2 s 18538 8500 18538 8500 4 fifo\[5\]\[3\]
rlabel metal1 s 19274 17612 19274 17612 4 fifo\[5\]\[4\]
rlabel metal1 s 24196 17646 24196 17646 4 fifo\[5\]\[5\]
rlabel metal1 s 28382 26860 28382 26860 4 fifo\[5\]\[6\]
rlabel metal1 s 27554 23290 27554 23290 4 fifo\[5\]\[7\]
rlabel metal2 s 30129 13294 30129 13294 4 fifo\[6\]\[0\]
rlabel metal1 s 30498 10030 30498 10030 4 fifo\[6\]\[1\]
rlabel metal2 s 24794 9214 24794 9214 4 fifo\[6\]\[2\]
rlabel metal1 s 20516 10030 20516 10030 4 fifo\[6\]\[3\]
rlabel metal2 s 27553 19346 27553 19346 4 fifo\[6\]\[4\]
rlabel metal2 s 29394 17510 29394 17510 4 fifo\[6\]\[5\]
rlabel metal1 s 30268 24038 30268 24038 4 fifo\[6\]\[6\]
rlabel metal1 s 29624 21114 29624 21114 4 fifo\[6\]\[7\]
rlabel metal1 s 12880 14042 12880 14042 4 fifo\[7\]\[0\]
rlabel metal1 s 14076 5338 14076 5338 4 fifo\[7\]\[1\]
rlabel metal1 s 8464 4250 8464 4250 4 fifo\[7\]\[2\]
rlabel metal1 s 8832 4726 8832 4726 4 fifo\[7\]\[3\]
rlabel metal1 s 12696 19482 12696 19482 4 fifo\[7\]\[4\]
rlabel metal2 s 7866 15028 7866 15028 4 fifo\[7\]\[5\]
rlabel metal1 s 8832 26418 8832 26418 4 fifo\[7\]\[6\]
rlabel metal1 s 8970 19890 8970 19890 4 fifo\[7\]\[7\]
rlabel metal1 s 25668 13906 25668 13906 4 fifo\[8\]\[0\]
rlabel metal1 s 27140 11730 27140 11730 4 fifo\[8\]\[1\]
rlabel metal1 s 23368 11730 23368 11730 4 fifo\[8\]\[2\]
rlabel metal1 s 20562 11186 20562 11186 4 fifo\[8\]\[3\]
rlabel metal1 s 21896 19482 21896 19482 4 fifo\[8\]\[4\]
rlabel metal2 s 27646 15164 27646 15164 4 fifo\[8\]\[5\]
rlabel metal1 s 25852 25330 25852 25330 4 fifo\[8\]\[6\]
rlabel metal1 s 25484 20910 25484 20910 4 fifo\[8\]\[7\]
rlabel metal2 s 21022 14586 21022 14586 4 fifo\[9\]\[0\]
rlabel metal1 s 26174 6222 26174 6222 4 fifo\[9\]\[1\]
rlabel metal1 s 22310 5202 22310 5202 4 fifo\[9\]\[2\]
rlabel metal1 s 19412 5678 19412 5678 4 fifo\[9\]\[3\]
rlabel metal1 s 20700 18938 20700 18938 4 fifo\[9\]\[4\]
rlabel metal2 s 23598 16626 23598 16626 4 fifo\[9\]\[5\]
rlabel metal1 s 24426 24854 24426 24854 4 fifo\[9\]\[6\]
rlabel metal1 s 24426 21590 24426 21590 4 fifo\[9\]\[7\]
rlabel metal2 s 17434 1520 17434 1520 4 full
rlabel metal2 s 20470 28458 20470 28458 4 head\[0\]
rlabel metal1 s 20056 31790 20056 31790 4 head\[1\]
rlabel metal1 s 19182 30702 19182 30702 4 head\[2\]
rlabel metal1 s 18676 27914 18676 27914 4 head\[3\]
rlabel metal1 s 12742 30838 12742 30838 4 head\[4\]
rlabel metal2 s 1702 20573 1702 20573 4 net1
rlabel metal1 s 7038 32266 7038 32266 4 net10
rlabel metal1 s 12696 18394 12696 18394 4 net100
rlabel metal1 s 20700 7786 20700 7786 4 net101
rlabel metal1 s 8418 26010 8418 26010 4 net102
rlabel metal2 s 30498 9792 30498 9792 4 net103
rlabel metal1 s 11960 14042 11960 14042 4 net104
rlabel metal1 s 8694 22746 8694 22746 4 net105
rlabel metal1 s 4094 14042 4094 14042 4 net106
rlabel metal1 s 27646 18258 27646 18258 4 net107
rlabel metal1 s 24610 16422 24610 16422 4 net108
rlabel metal1 s 3680 14994 3680 14994 4 net109
rlabel metal2 s 18952 15130 18952 15130 4 net11
rlabel metal1 s 25760 6290 25760 6290 4 net110
rlabel metal1 s 20240 18258 20240 18258 4 net111
rlabel metal1 s 29072 22610 29072 22610 4 net112
rlabel metal1 s 17848 6290 17848 6290 4 net113
rlabel metal1 s 7268 18666 7268 18666 4 net114
rlabel metal1 s 8648 9962 8648 9962 4 net115
rlabel metal1 s 17572 8874 17572 8874 4 net116
rlabel metal1 s 26726 25874 26726 25874 4 net117
rlabel metal1 s 27462 27098 27462 27098 4 net118
rlabel metal1 s 9292 20570 9292 20570 4 net119
rlabel metal1 s 20654 2414 20654 2414 4 net12
rlabel metal1 s 10672 8602 10672 8602 4 net120
rlabel metal2 s 6946 11424 6946 11424 4 net121
rlabel metal1 s 19918 12138 19918 12138 4 net122
rlabel metal1 s 24978 17306 24978 17306 4 net123
rlabel metal1 s 4370 11866 4370 11866 4 net124
rlabel metal1 s 22080 19754 22080 19754 4 net125
rlabel metal1 s 4600 10642 4600 10642 4 net126
rlabel metal1 s 6072 25194 6072 25194 4 net127
rlabel metal1 s 4416 11050 4416 11050 4 net128
rlabel metal1 s 24058 27098 24058 27098 4 net129
rlabel metal1 s 4347 2414 4347 2414 4 net13
rlabel metal1 s 25070 25194 25070 25194 4 net130
rlabel metal1 s 9108 5202 9108 5202 4 net131
rlabel metal1 s 18768 8466 18768 8466 4 net132
rlabel metal2 s 6762 26384 6762 26384 4 net133
rlabel metal1 s 10396 6630 10396 6630 4 net134
rlabel metal1 s 25024 9962 25024 9962 4 net135
rlabel metal1 s 5566 21114 5566 21114 4 net136
rlabel metal1 s 6716 15130 6716 15130 4 net137
rlabel metal1 s 4508 19754 4508 19754 4 net138
rlabel metal1 s 27738 26350 27738 26350 4 net139
rlabel metal1 s 8464 2346 8464 2346 4 net14
rlabel metal1 s 9660 10778 9660 10778 4 net140
rlabel metal1 s 14720 5610 14720 5610 4 net141
rlabel metal2 s 27370 13328 27370 13328 4 net142
rlabel metal1 s 29946 24854 29946 24854 4 net143
rlabel metal1 s 6302 11866 6302 11866 4 net144
rlabel metal1 s 7360 7786 7360 7786 4 net145
rlabel metal1 s 7820 7378 7820 7378 4 net146
rlabel metal1 s 4416 9962 4416 9962 4 net147
rlabel metal1 s 9476 28050 9476 28050 4 net148
rlabel metal1 s 5244 25874 5244 25874 4 net149
rlabel metal1 s 2277 12886 2277 12886 4 net15
rlabel metal1 s 6670 21658 6670 21658 4 net150
rlabel metal1 s 18722 13498 18722 13498 4 net151
rlabel metal1 s 15272 7378 15272 7378 4 net152
rlabel metal1 s 8510 4794 8510 4794 4 net153
rlabel metal1 s 11270 28050 11270 28050 4 net154
rlabel metal1 s 7222 5678 7222 5678 4 net155
rlabel metal1 s 12190 31314 12190 31314 4 net156
rlabel metal1 s 6670 7514 6670 7514 4 net157
rlabel metal1 s 16836 30226 16836 30226 4 net158
rlabel metal1 s 11224 4182 11224 4182 4 net159
rlabel metal2 s 15042 4352 15042 4352 4 net16
rlabel metal1 s 17986 31382 17986 31382 4 net160
rlabel metal1 s 18032 30906 18032 30906 4 net161
rlabel metal1 s 10304 4250 10304 4250 4 net162
rlabel metal1 s 23552 23630 23552 23630 4 net163
rlabel metal1 s 23322 24174 23322 24174 4 net164
rlabel metal1 s 29256 23698 29256 23698 4 net165
rlabel metal1 s 28290 22610 28290 22610 4 net166
rlabel metal1 s 12006 3366 12006 3366 4 net17
rlabel metal1 s 22080 20400 22080 20400 4 net18
rlabel metal3 s 10718 24667 10718 24667 4 net19
rlabel metal1 s 29348 2618 29348 2618 4 net2
rlabel metal2 s 13570 31586 13570 31586 4 net20
rlabel metal2 s 24702 31926 24702 31926 4 net21
rlabel metal1 s 17342 2414 17342 2414 4 net22
rlabel metal2 s 14400 8466 14400 8466 4 net23
rlabel metal1 s 25622 24718 25622 24718 4 net24
rlabel metal1 s 25162 24072 25162 24072 4 net25
rlabel metal1 s 21827 10030 21827 10030 4 net26
rlabel metal1 s 21111 10030 21111 10030 4 net27
rlabel metal1 s 15732 14042 15732 14042 4 net28
rlabel metal1 s 12098 24922 12098 24922 4 net29
rlabel metal1 s 16698 6664 16698 6664 4 net3
rlabel metal1 s 15088 17578 15088 17578 4 net30
rlabel metal1 s 15088 8942 15088 8942 4 net31
rlabel metal1 s 11040 20910 11040 20910 4 net32
rlabel metal1 s 11132 16218 11132 16218 4 net33
rlabel metal1 s 13478 17306 13478 17306 4 net34
rlabel metal1 s 14720 13226 14720 13226 4 net35
rlabel metal1 s 8464 18258 8464 18258 4 net36
rlabel metal1 s 19136 18394 19136 18394 4 net37
rlabel metal1 s 21804 18666 21804 18666 4 net38
rlabel metal1 s 19918 19482 19918 19482 4 net39
rlabel metal1 s 8418 7514 8418 7514 4 net4
rlabel metal1 s 25024 21658 25024 21658 4 net40
rlabel metal1 s 4416 18666 4416 18666 4 net41
rlabel metal2 s 13018 9146 13018 9146 4 net42
rlabel metal2 s 29578 21760 29578 21760 4 net43
rlabel metal1 s 13386 14382 13386 14382 4 net44
rlabel metal1 s 21390 14042 21390 14042 4 net45
rlabel metal1 s 12144 10778 12144 10778 4 net46
rlabel metal1 s 25438 20570 25438 20570 4 net47
rlabel metal1 s 15870 18394 15870 18394 4 net48
rlabel metal1 s 23092 15402 23092 15402 4 net49
rlabel metal2 s 13478 18938 13478 18938 4 net5
rlabel metal1 s 14352 14042 14352 14042 4 net50
rlabel metal1 s 22678 15130 22678 15130 4 net51
rlabel metal1 s 13616 19346 13616 19346 4 net52
rlabel metal1 s 11316 18734 11316 18734 4 net53
rlabel metal2 s 27922 20706 27922 20706 4 net54
rlabel metal1 s 27600 16082 27600 16082 4 net55
rlabel metal1 s 25162 12954 25162 12954 4 net56
rlabel metal1 s 22218 11118 22218 11118 4 net57
rlabel metal1 s 25024 6698 25024 6698 4 net58
rlabel metal1 s 16192 12138 16192 12138 4 net59
rlabel metal1 s 15226 16048 15226 16048 4 net6
rlabel metal1 s 30038 12138 30038 12138 4 net60
rlabel metal1 s 24150 25262 24150 25262 4 net61
rlabel metal1 s 25208 22746 25208 22746 4 net62
rlabel metal1 s 7820 16558 7820 16558 4 net63
rlabel metal1 s 8694 24922 8694 24922 4 net64
rlabel metal1 s 18170 14246 18170 14246 4 net65
rlabel metal2 s 29026 21114 29026 21114 4 net66
rlabel metal1 s 20792 9146 20792 9146 4 net67
rlabel metal1 s 28612 17306 28612 17306 4 net68
rlabel metal1 s 30176 17306 30176 17306 4 net69
rlabel metal1 s 5796 25942 5796 25942 4 net7
rlabel metal1 s 8602 19482 8602 19482 4 net70
rlabel metal1 s 10212 27098 10212 27098 4 net71
rlabel metal2 s 4646 16354 4646 16354 4 net72
rlabel metal1 s 26266 15334 26266 15334 4 net73
rlabel metal1 s 19964 9962 19964 9962 4 net74
rlabel metal1 s 29256 13906 29256 13906 4 net75
rlabel metal1 s 12604 6290 12604 6290 4 net76
rlabel metal1 s 18998 5610 18998 5610 4 net77
rlabel metal2 s 29026 24344 29026 24344 4 net78
rlabel metal1 s 26312 10778 26312 10778 4 net79
rlabel metal1 s 8142 21658 8142 21658 4 net8
rlabel metal1 s 27416 18394 27416 18394 4 net80
rlabel metal1 s 22586 7786 22586 7786 4 net81
rlabel metal1 s 27508 7378 27508 7378 4 net82
rlabel metal1 s 20792 5678 20792 5678 4 net83
rlabel metal1 s 25024 8874 25024 8874 4 net84
rlabel metal1 s 27416 21998 27416 21998 4 net85
rlabel metal1 s 14720 7786 14720 7786 4 net86
rlabel metal1 s 19642 14484 19642 14484 4 net87
rlabel metal1 s 15088 10778 15088 10778 4 net88
rlabel metal2 s 23322 12410 23322 12410 4 net89
rlabel metal2 s 3818 24276 3818 24276 4 net9
rlabel metal1 s 21804 5338 21804 5338 4 net90
rlabel metal1 s 27692 8466 27692 8466 4 net91
rlabel metal2 s 5474 22848 5474 22848 4 net92
rlabel metal1 s 5336 17306 5336 17306 4 net93
rlabel metal1 s 28612 9622 28612 9622 4 net94
rlabel metal1 s 19872 11050 19872 11050 4 net95
rlabel metal1 s 18170 18734 18170 18734 4 net96
rlabel metal1 s 27784 10778 27784 10778 4 net97
rlabel metal1 s 9844 15130 9844 15130 4 net98
rlabel metal2 s 7958 14790 7958 14790 4 net99
rlabel metal3 s 820 24548 820 24548 4 pop
rlabel metal1 s 1380 32402 1380 32402 4 push
rlabel metal2 s 31510 13753 31510 13753 4 rst
rlabel metal2 s 20562 25602 20562 25602 4 tail\[0\]
rlabel metal2 s 20470 24225 20470 24225 4 tail\[1\]
rlabel metal2 s 19918 26180 19918 26180 4 tail\[2\]
rlabel metal1 s 20194 24174 20194 24174 4 tail\[3\]
rlabel metal1 s 12144 28730 12144 28730 4 tail\[4\]
flabel metal5 s 1056 30046 31880 30446 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 24046 31880 24446 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 18046 31880 18446 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 12046 31880 12446 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 6046 31880 6446 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal4 s 28908 2128 29308 32688 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 22908 2128 23308 32688 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 16908 2128 17308 32688 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 10908 2128 11308 32688 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 4908 2128 5308 32688 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal5 s 1056 29306 31880 29706 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 23306 31880 23706 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 17306 31880 17706 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 11306 31880 11706 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 5306 31880 5706 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal4 s 28168 2128 28568 32688 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 22168 2128 22568 32688 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 16168 2128 16568 32688 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 10168 2128 10568 32688 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 4168 2128 4568 32688 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal3 s 32174 31968 32974 32088 0 FreeSans 600 0 0 0 clk
port 3 nsew
flabel metal3 s 0 30608 800 30728 0 FreeSans 600 0 0 0 data_in[0]
port 4 nsew
flabel metal2 s 28998 0 29054 800 0 FreeSans 280 90 0 0 data_in[1]
port 5 nsew
flabel metal3 s 0 6128 800 6248 0 FreeSans 600 0 0 0 data_in[2]
port 6 nsew
flabel metal3 s 0 18368 800 18488 0 FreeSans 600 0 0 0 data_in[3]
port 7 nsew
flabel metal2 s 7102 34318 7158 35118 0 FreeSans 280 90 0 0 data_in[4]
port 8 nsew
flabel metal2 s 12898 34318 12954 35118 0 FreeSans 280 90 0 0 data_in[5]
port 9 nsew
flabel metal2 s 30286 34318 30342 35118 0 FreeSans 280 90 0 0 data_in[6]
port 10 nsew
flabel metal3 s 32174 7488 32974 7608 0 FreeSans 600 0 0 0 data_in[7]
port 11 nsew
flabel metal2 s 23202 0 23258 800 0 FreeSans 280 90 0 0 data_out[0]
port 12 nsew
flabel metal2 s 18 0 74 800 0 FreeSans 280 90 0 0 data_out[1]
port 13 nsew
flabel metal2 s 5814 0 5870 800 0 FreeSans 280 90 0 0 data_out[2]
port 14 nsew
flabel metal3 s 0 12248 800 12368 0 FreeSans 600 0 0 0 data_out[3]
port 15 nsew
flabel metal3 s 32174 1368 32974 1488 0 FreeSans 600 0 0 0 data_out[4]
port 16 nsew
flabel metal2 s 11610 0 11666 800 0 FreeSans 280 90 0 0 data_out[5]
port 17 nsew
flabel metal3 s 32174 19728 32974 19848 0 FreeSans 600 0 0 0 data_out[6]
port 18 nsew
flabel metal3 s 32174 25848 32974 25968 0 FreeSans 600 0 0 0 data_out[7]
port 19 nsew
flabel metal2 s 18694 34318 18750 35118 0 FreeSans 280 90 0 0 empty
port 20 nsew
flabel metal2 s 24490 34318 24546 35118 0 FreeSans 280 90 0 0 error
port 21 nsew
flabel metal2 s 17406 0 17462 800 0 FreeSans 280 90 0 0 full
port 22 nsew
flabel metal3 s 0 24488 800 24608 0 FreeSans 600 0 0 0 pop
port 23 nsew
flabel metal2 s 1306 34318 1362 35118 0 FreeSans 280 90 0 0 push
port 24 nsew
flabel metal3 s 32174 13608 32974 13728 0 FreeSans 600 0 0 0 rst
port 25 nsew
<< properties >>
string FIXED_BBOX 0 0 32974 35118
<< end >>
