* NGSPICE file created from fifo.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

.subckt fifo VGND VPWR clk data_in[0] data_in[1] data_in[2] data_in[3] data_in[4]
+ data_in[5] data_in[6] data_in[7] data_out[0] data_out[1] data_out[2] data_out[3]
+ data_out[4] data_out[5] data_out[6] data_out[7] empty error full pop push rst
XTAP_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0985_ clknet_4_2_0_clk _0025_ _0006_ VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_196 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0770_ _0372_ VGND VGND VPWR VPWR _0072_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_4_12_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_12_0_clk sky130_fd_sc_hd__clkbuf_8
X_0968_ net145 net3 _0480_ VGND VGND VPWR VPWR _0483_ sky130_fd_sc_hd__mux2_1
X_0899_ _0444_ VGND VGND VPWR VPWR _0129_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0822_ _0401_ VGND VGND VPWR VPWR _0095_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0753_ _0362_ VGND VGND VPWR VPWR _0065_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0684_ net28 _0315_ _0320_ VGND VGND VPWR VPWR _0321_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1098_ clknet_4_2_0_clk _0137_ VGND VGND VPWR VPWR fifo\[12\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1021_ clknet_4_15_0_clk _0060_ VGND VGND VPWR VPWR fifo\[2\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_0805_ net84 _0324_ _0389_ VGND VGND VPWR VPWR _0392_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0667_ _0314_ VGND VGND VPWR VPWR _0009_ sky130_fd_sc_hd__inv_2
X_0598_ _0262_ VGND VGND VPWR VPWR _0025_ sky130_fd_sc_hd__clkbuf_1
X_0736_ net107 _0328_ _0348_ VGND VGND VPWR VPWR _0353_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold63 fifo\[9\]\[2\] VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 fifo\[14\]\[2\] VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__dlygate4sd3_1
Xhold30 fifo\[8\]\[2\] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 fifo\[8\]\[1\] VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 fifo\[6\]\[5\] VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 fifo\[14\]\[7\] VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__dlygate4sd3_1
Xhold96 fifo\[5\]\[5\] VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0521_ head\[2\] _0191_ _0190_ VGND VGND VPWR VPWR _0194_ sky130_fd_sc_hd__and3_1
XTAP_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1004_ clknet_4_4_0_clk _0043_ VGND VGND VPWR VPWR fifo\[0\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0719_ net55 _0330_ _0337_ VGND VGND VPWR VPWR _0343_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_204 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput20 net20 VGND VGND VPWR VPWR empty sky130_fd_sc_hd__clkbuf_4
XFILLER_0_53_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0504_ _0179_ _0180_ VGND VGND VPWR VPWR _0181_ sky130_fd_sc_hd__nand2_1
XTAP_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0984_ clknet_4_1_0_clk _0024_ _0005_ VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_60 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0967_ _0482_ VGND VGND VPWR VPWR _0159_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0898_ net128 net4 _0440_ VGND VGND VPWR VPWR _0444_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0821_ net141 _0322_ _0399_ VGND VGND VPWR VPWR _0401_ sky130_fd_sc_hd__mux2_1
X_0752_ net134 _0326_ _0358_ VGND VGND VPWR VPWR _0362_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0683_ _0319_ VGND VGND VPWR VPWR _0320_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1097_ clknet_4_8_0_clk _0136_ VGND VGND VPWR VPWR fifo\[12\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_118 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_4_11_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_11_0_clk sky130_fd_sc_hd__clkbuf_8
X_1020_ clknet_4_11_0_clk _0059_ VGND VGND VPWR VPWR fifo\[2\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0804_ _0391_ VGND VGND VPWR VPWR _0087_ sky130_fd_sc_hd__clkbuf_1
X_0735_ _0352_ VGND VGND VPWR VPWR _0057_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0666_ _0314_ VGND VGND VPWR VPWR _0008_ sky130_fd_sc_hd__inv_2
X_0597_ net16 _0261_ _0172_ VGND VGND VPWR VPWR _0262_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_243 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_151 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold75 fifo\[7\]\[6\] VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__dlygate4sd3_1
Xhold20 fifo\[8\]\[7\] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 fifo\[6\]\[4\] VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 fifo\[12\]\[3\] VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 fifo\[12\]\[1\] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 fifo\[14\]\[1\] VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 fifo\[13\]\[3\] VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 fifo\[2\]\[5\] VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0520_ _0191_ _0192_ VGND VGND VPWR VPWR _0193_ sky130_fd_sc_hd__and2_1
XTAP_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1003_ clknet_4_6_0_clk _0042_ VGND VGND VPWR VPWR fifo\[0\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_0718_ _0342_ VGND VGND VPWR VPWR _0050_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0649_ net12 _0309_ _0172_ VGND VGND VPWR VPWR _0310_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_216 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput21 net21 VGND VGND VPWR VPWR error sky130_fd_sc_hd__clkbuf_4
XFILLER_0_53_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0503_ tail\[0\] VGND VGND VPWR VPWR _0180_ sky130_fd_sc_hd__buf_2
XTAP_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0983_ clknet_4_0_0_clk _0023_ _0004_ VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0966_ net86 net2 _0480_ VGND VGND VPWR VPWR _0482_ sky130_fd_sc_hd__mux2_1
X_0897_ _0443_ VGND VGND VPWR VPWR _0128_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0751_ _0361_ VGND VGND VPWR VPWR _0064_ sky130_fd_sc_hd__clkbuf_1
X_0820_ _0400_ VGND VGND VPWR VPWR _0094_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0682_ _0196_ _0316_ _0317_ _0318_ VGND VGND VPWR VPWR _0319_ sky130_fd_sc_hd__and4b_1
X_1096_ clknet_4_10_0_clk _0135_ VGND VGND VPWR VPWR fifo\[12\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0949_ _0472_ VGND VGND VPWR VPWR _0151_ sky130_fd_sc_hd__clkbuf_1
X_0665_ _0314_ VGND VGND VPWR VPWR _0007_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0734_ net67 _0326_ _0348_ VGND VGND VPWR VPWR _0352_ sky130_fd_sc_hd__mux2_1
X_0803_ net94 _0322_ _0389_ VGND VGND VPWR VPWR _0391_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0596_ _0255_ _0257_ _0259_ _0260_ VGND VGND VPWR VPWR _0261_ sky130_fd_sc_hd__o31a_1
XFILLER_0_47_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1079_ clknet_4_1_0_clk _0118_ VGND VGND VPWR VPWR fifo\[10\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_255 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold65 fifo\[13\]\[7\] VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 fifo\[1\]\[4\] VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 fifo\[7\]\[7\] VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__dlygate4sd3_1
Xhold10 fifo\[14\]\[4\] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 fifo\[4\]\[4\] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 fifo\[5\]\[2\] VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 fifo\[2\]\[1\] VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 fifo\[4\]\[0\] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 fifo\[10\]\[7\] VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1002_ clknet_4_0_0_clk _0041_ VGND VGND VPWR VPWR fifo\[0\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0717_ net125 _0328_ _0337_ VGND VGND VPWR VPWR _0342_ sky130_fd_sc_hd__mux2_1
X_0648_ _0303_ _0305_ _0307_ _0308_ VGND VGND VPWR VPWR _0309_ sky130_fd_sc_hd__o31a_1
X_0579_ fifo\[4\]\[5\] _0212_ _0244_ VGND VGND VPWR VPWR _0245_ sky130_fd_sc_hd__a21o_1
XFILLER_0_50_228 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_4_10_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_10_0_clk sky130_fd_sc_hd__clkbuf_8
Xoutput22 net22 VGND VGND VPWR VPWR full sky130_fd_sc_hd__clkbuf_4
XFILLER_0_9_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0502_ tail\[1\] VGND VGND VPWR VPWR _0179_ sky130_fd_sc_hd__buf_2
XTAP_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0982_ clknet_4_2_0_clk _0022_ _0003_ VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0896_ net147 net3 _0440_ VGND VGND VPWR VPWR _0443_ sky130_fd_sc_hd__mux2_1
X_0965_ _0481_ VGND VGND VPWR VPWR _0158_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0681_ head\[3\] head\[2\] VGND VGND VPWR VPWR _0318_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0750_ net120 _0324_ _0358_ VGND VGND VPWR VPWR _0361_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1095_ clknet_4_9_0_clk _0134_ VGND VGND VPWR VPWR fifo\[12\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0948_ net91 net2 _0470_ VGND VGND VPWR VPWR _0472_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0879_ _0433_ VGND VGND VPWR VPWR _0120_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0802_ _0390_ VGND VGND VPWR VPWR _0086_ sky130_fd_sc_hd__clkbuf_1
X_0664_ _0314_ VGND VGND VPWR VPWR _0006_ sky130_fd_sc_hd__inv_2
X_0733_ _0351_ VGND VGND VPWR VPWR _0056_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0595_ fifo\[0\]\[4\] _0223_ VGND VGND VPWR VPWR _0260_ sky130_fd_sc_hd__or2_1
X_1078_ clknet_4_13_0_clk _0117_ VGND VGND VPWR VPWR fifo\[9\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold11 fifo\[8\]\[4\] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 fifo\[12\]\[5\] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 fifo\[3\]\[6\] VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 fifo\[5\]\[1\] VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 fifo\[4\]\[2\] VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 fifo\[13\]\[2\] VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 fifo\[2\]\[0\] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 fifo\[10\]\[0\] VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 fifo\[13\]\[5\] VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1001_ clknet_4_2_0_clk _0040_ VGND VGND VPWR VPWR fifo\[0\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0716_ _0341_ VGND VGND VPWR VPWR _0049_ sky130_fd_sc_hd__clkbuf_1
X_0647_ fifo\[0\]\[0\] _0223_ VGND VGND VPWR VPWR _0308_ sky130_fd_sc_hd__or2_1
X_0578_ fifo\[11\]\[5\] _0213_ _0214_ fifo\[13\]\[5\] VGND VGND VPWR VPWR _0244_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_204 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput12 net12 VGND VGND VPWR VPWR data_out[0] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0501_ _0170_ _0171_ net9 VGND VGND VPWR VPWR _0178_ sky130_fd_sc_hd__a21bo_1
XTAP_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0981_ clknet_4_2_0_clk _0021_ _0002_ VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold130 fifo\[15\]\[3\] VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0964_ net44 net1 _0480_ VGND VGND VPWR VPWR _0481_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0895_ _0442_ VGND VGND VPWR VPWR _0127_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0680_ head\[1\] _0313_ VGND VGND VPWR VPWR _0317_ sky130_fd_sc_hd__nor2_2
XFILLER_0_36_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1094_ clknet_4_5_0_clk _0133_ VGND VGND VPWR VPWR fifo\[11\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0947_ _0471_ VGND VGND VPWR VPWR _0150_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0878_ net155 net3 _0430_ VGND VGND VPWR VPWR _0433_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0801_ net75 _0315_ _0389_ VGND VGND VPWR VPWR _0390_ sky130_fd_sc_hd__mux2_1
X_0732_ net135 _0324_ _0348_ VGND VGND VPWR VPWR _0351_ sky130_fd_sc_hd__mux2_1
X_0663_ _0314_ VGND VGND VPWR VPWR _0005_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0594_ fifo\[3\]\[4\] net23 _0219_ fifo\[15\]\[4\] _0258_ VGND VGND VPWR VPWR _0259_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1077_ clknet_4_15_0_clk _0116_ VGND VGND VPWR VPWR fifo\[9\]\[6\] sky130_fd_sc_hd__dfxtp_1
Xhold34 fifo\[9\]\[6\] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__dlygate4sd3_1
Xhold12 fifo\[9\]\[4\] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 fifo\[12\]\[2\] VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 fifo\[7\]\[0\] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 fifo\[11\]\[5\] VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 fifo\[4\]\[7\] VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 fifo\[14\]\[3\] VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 fifo\[6\]\[1\] VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1000_ clknet_4_3_0_clk _0039_ VGND VGND VPWR VPWR fifo\[0\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0715_ net122 _0326_ _0337_ VGND VGND VPWR VPWR _0341_ sky130_fd_sc_hd__mux2_1
X_0646_ fifo\[3\]\[0\] net23 _0219_ fifo\[15\]\[0\] _0306_ VGND VGND VPWR VPWR _0307_
+ sky130_fd_sc_hd__a221o_1
X_0577_ _0239_ _0240_ _0241_ _0242_ VGND VGND VPWR VPWR _0243_ sky130_fd_sc_hd__or4_1
XFILLER_0_25_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput13 net13 VGND VGND VPWR VPWR data_out[1] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0500_ _0176_ VGND VGND VPWR VPWR _0177_ sky130_fd_sc_hd__inv_2
XTAP_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_274 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_110 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0629_ _0287_ _0288_ _0289_ _0290_ VGND VGND VPWR VPWR _0291_ sky130_fd_sc_hd__or4_1
XFILLER_0_31_241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0980_ clknet_4_7_0_clk _0020_ _0001_ VGND VGND VPWR VPWR tail\[4\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_38_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold131 head\[3\] VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold120 fifo\[11\]\[2\] VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_160 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0963_ _0479_ VGND VGND VPWR VPWR _0480_ sky130_fd_sc_hd__buf_4
XFILLER_0_39_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0894_ net121 net2 _0440_ VGND VGND VPWR VPWR _0442_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1093_ clknet_4_5_0_clk _0132_ VGND VGND VPWR VPWR fifo\[11\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0877_ _0432_ VGND VGND VPWR VPWR _0119_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_314 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0946_ net65 net1 _0470_ VGND VGND VPWR VPWR _0471_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_196 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_174 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0800_ _0388_ VGND VGND VPWR VPWR _0389_ sky130_fd_sc_hd__buf_4
XFILLER_0_12_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0731_ _0350_ VGND VGND VPWR VPWR _0055_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_67 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0662_ _0314_ VGND VGND VPWR VPWR _0004_ sky130_fd_sc_hd__inv_2
X_0593_ fifo\[7\]\[4\] _0175_ _0220_ fifo\[10\]\[4\] VGND VGND VPWR VPWR _0258_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1076_ clknet_4_9_0_clk _0115_ VGND VGND VPWR VPWR fifo\[9\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0929_ _0461_ VGND VGND VPWR VPWR _0142_ sky130_fd_sc_hd__clkbuf_1
Xhold35 fifo\[12\]\[7\] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__dlygate4sd3_1
Xhold13 fifo\[9\]\[7\] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__dlygate4sd3_1
Xhold57 fifo\[6\]\[2\] VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 fifo\[8\]\[3\] VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 fifo\[13\]\[0\] VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 fifo\[8\]\[5\] VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 fifo\[9\]\[5\] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0645_ fifo\[7\]\[0\] _0175_ _0220_ fifo\[10\]\[0\] VGND VGND VPWR VPWR _0306_ sky130_fd_sc_hd__a22o_1
X_0714_ _0340_ VGND VGND VPWR VPWR _0048_ sky130_fd_sc_hd__clkbuf_1
X_0576_ fifo\[9\]\[5\] _0208_ _0209_ fifo\[12\]\[5\] VGND VGND VPWR VPWR _0242_ sky130_fd_sc_hd__a22o_1
X_1059_ clknet_4_6_0_clk _0098_ VGND VGND VPWR VPWR fifo\[7\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput14 net14 VGND VGND VPWR VPWR data_out[2] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_34_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0628_ fifo\[9\]\[1\] _0208_ _0209_ fifo\[12\]\[1\] VGND VGND VPWR VPWR _0290_ sky130_fd_sc_hd__a22o_1
X_0559_ _0226_ VGND VGND VPWR VPWR _0028_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold110 fifo\[10\]\[5\] VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__dlygate4sd3_1
Xhold121 fifo\[15\]\[6\] VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__dlygate4sd3_1
Xhold132 net17 VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_172 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0962_ _0001_ _0191_ _0189_ _0192_ VGND VGND VPWR VPWR _0479_ sky130_fd_sc_hd__and4_1
XFILLER_0_40_55 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_228 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0893_ _0441_ VGND VGND VPWR VPWR _0126_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1092_ clknet_4_4_0_clk _0131_ VGND VGND VPWR VPWR fifo\[11\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_0945_ _0469_ VGND VGND VPWR VPWR _0470_ sky130_fd_sc_hd__buf_4
XFILLER_0_42_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0876_ net76 net2 _0430_ VGND VGND VPWR VPWR _0432_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0661_ _0314_ VGND VGND VPWR VPWR _0003_ sky130_fd_sc_hd__inv_2
X_0730_ net103 _0322_ _0348_ VGND VGND VPWR VPWR _0350_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_79 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0592_ fifo\[4\]\[4\] _0212_ _0256_ VGND VGND VPWR VPWR _0257_ sky130_fd_sc_hd__a21o_1
X_1075_ clknet_4_12_0_clk _0114_ VGND VGND VPWR VPWR fifo\[9\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0859_ _0422_ VGND VGND VPWR VPWR _0111_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0928_ net106 net1 _0460_ VGND VGND VPWR VPWR _0461_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold58 fifo\[5\]\[7\] VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 fifo\[12\]\[4\] VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 fifo\[15\]\[4\] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 fifo\[6\]\[3\] VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 fifo\[15\]\[5\] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__dlygate4sd3_1
Xhold14 fifo\[13\]\[4\] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0713_ net89 _0324_ _0337_ VGND VGND VPWR VPWR _0340_ sky130_fd_sc_hd__mux2_1
X_0644_ fifo\[4\]\[0\] _0212_ _0304_ VGND VGND VPWR VPWR _0305_ sky130_fd_sc_hd__a21o_1
X_0575_ fifo\[14\]\[5\] _0205_ _0206_ fifo\[5\]\[5\] VGND VGND VPWR VPWR _0241_ sky130_fd_sc_hd__a22o_1
X_1058_ clknet_4_0_0_clk _0097_ VGND VGND VPWR VPWR fifo\[7\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput15 net15 VGND VGND VPWR VPWR data_out[3] sky130_fd_sc_hd__clkbuf_4
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0558_ net19 _0225_ _0172_ VGND VGND VPWR VPWR _0226_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_88 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0627_ fifo\[14\]\[1\] _0205_ _0206_ fifo\[5\]\[1\] VGND VGND VPWR VPWR _0289_ sky130_fd_sc_hd__a22o_1
X_0489_ tail\[2\] head\[2\] VGND VGND VPWR VPWR _0166_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_48_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold133 head\[1\] VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__dlygate4sd3_1
Xhold122 fifo\[13\]\[6\] VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__dlygate4sd3_1
Xhold100 fifo\[11\]\[6\] VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__dlygate4sd3_1
Xhold111 fifo\[11\]\[4\] VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_51_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0961_ _0478_ VGND VGND VPWR VPWR _0157_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0892_ net109 net1 _0440_ VGND VGND VPWR VPWR _0441_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1091_ clknet_4_4_0_clk _0130_ VGND VGND VPWR VPWR fifo\[11\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0944_ _0196_ _0316_ _0192_ _0346_ VGND VGND VPWR VPWR _0469_ sky130_fd_sc_hd__and4b_1
XFILLER_0_27_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0875_ _0431_ VGND VGND VPWR VPWR _0118_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0660_ _0314_ VGND VGND VPWR VPWR _0002_ sky130_fd_sc_hd__inv_2
X_0591_ fifo\[11\]\[4\] _0213_ _0214_ fifo\[13\]\[4\] VGND VGND VPWR VPWR _0256_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1074_ clknet_4_8_0_clk _0113_ VGND VGND VPWR VPWR fifo\[9\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0927_ _0459_ VGND VGND VPWR VPWR _0460_ sky130_fd_sc_hd__clkbuf_4
X_0858_ net110 _0322_ _0420_ VGND VGND VPWR VPWR _0422_ sky130_fd_sc_hd__mux2_1
X_0789_ net132 _0326_ _0379_ VGND VGND VPWR VPWR _0383_ sky130_fd_sc_hd__mux2_1
Xhold37 fifo\[4\]\[6\] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 fifo\[10\]\[4\] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 fifo\[15\]\[1\] VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__dlygate4sd3_1
Xhold15 fifo\[0\]\[2\] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__dlygate4sd3_1
Xhold48 fifo\[6\]\[0\] VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0712_ _0339_ VGND VGND VPWR VPWR _0047_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_171 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0643_ fifo\[11\]\[0\] _0213_ _0214_ fifo\[13\]\[0\] VGND VGND VPWR VPWR _0304_ sky130_fd_sc_hd__a22o_1
X_0574_ fifo\[1\]\[5\] net25 net24 fifo\[8\]\[5\] VGND VGND VPWR VPWR _0240_ sky130_fd_sc_hd__a22o_1
X_1126_ clknet_4_5_0_clk _0165_ VGND VGND VPWR VPWR fifo\[15\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_1057_ clknet_4_0_0_clk _0096_ VGND VGND VPWR VPWR fifo\[7\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput16 net16 VGND VGND VPWR VPWR data_out[4] sky130_fd_sc_hd__buf_2
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
X_0557_ _0211_ _0216_ _0222_ _0224_ VGND VGND VPWR VPWR _0225_ sky130_fd_sc_hd__o31a_1
X_0626_ fifo\[1\]\[1\] net25 net24 fifo\[8\]\[1\] VGND VGND VPWR VPWR _0288_ sky130_fd_sc_hd__a22o_1
X_1109_ clknet_4_5_0_clk _0148_ VGND VGND VPWR VPWR fifo\[13\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_116 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold134 head\[2\] VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__dlygate4sd3_1
Xhold112 fifo\[5\]\[6\] VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__dlygate4sd3_1
Xhold123 fifo\[15\]\[7\] VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__dlygate4sd3_1
Xhold101 fifo\[11\]\[3\] VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__dlygate4sd3_1
X_0609_ _0267_ _0269_ _0271_ _0272_ VGND VGND VPWR VPWR _0273_ sky130_fd_sc_hd__o31a_1
XFILLER_0_51_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0960_ net112 net8 _0470_ VGND VGND VPWR VPWR _0478_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0891_ _0439_ VGND VGND VPWR VPWR _0440_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1090_ clknet_4_1_0_clk _0129_ VGND VGND VPWR VPWR fifo\[11\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_0943_ _0468_ VGND VGND VPWR VPWR _0149_ sky130_fd_sc_hd__clkbuf_1
X_0874_ net104 net1 _0430_ VGND VGND VPWR VPWR _0431_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_111 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0590_ _0251_ _0252_ _0253_ _0254_ VGND VGND VPWR VPWR _0255_ sky130_fd_sc_hd__or4_1
X_1073_ clknet_4_8_0_clk _0112_ VGND VGND VPWR VPWR fifo\[9\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0926_ head\[0\] _0190_ _0192_ _0317_ VGND VGND VPWR VPWR _0459_ sky130_fd_sc_hd__and4_1
XFILLER_0_11_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0857_ _0421_ VGND VGND VPWR VPWR _0110_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold16 fifo\[6\]\[7\] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 fifo\[1\]\[7\] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__dlygate4sd3_1
X_0788_ _0382_ VGND VGND VPWR VPWR _0080_ sky130_fd_sc_hd__clkbuf_1
Xhold38 fifo\[14\]\[0\] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 fifo\[10\]\[1\] VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_220 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0711_ net97 _0322_ _0337_ VGND VGND VPWR VPWR _0339_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0642_ _0299_ _0300_ _0301_ _0302_ VGND VGND VPWR VPWR _0303_ sky130_fd_sc_hd__or4_1
X_0573_ fifo\[2\]\[5\] net27 _0199_ fifo\[6\]\[5\] net26 VGND VGND VPWR VPWR _0239_
+ sky130_fd_sc_hd__a221o_1
X_1125_ clknet_4_5_0_clk _0164_ VGND VGND VPWR VPWR fifo\[15\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1056_ clknet_4_2_0_clk _0095_ VGND VGND VPWR VPWR fifo\[7\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0909_ _0449_ VGND VGND VPWR VPWR _0450_ sky130_fd_sc_hd__buf_4
Xoutput17 net17 VGND VGND VPWR VPWR data_out[5] sky130_fd_sc_hd__clkbuf_4
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0625_ fifo\[2\]\[1\] net27 _0199_ fifo\[6\]\[1\] net26 VGND VGND VPWR VPWR _0287_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_25_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0556_ fifo\[0\]\[7\] _0223_ VGND VGND VPWR VPWR _0224_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_91 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1039_ clknet_4_9_0_clk _0078_ VGND VGND VPWR VPWR fifo\[5\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_1108_ clknet_4_4_0_clk _0147_ VGND VGND VPWR VPWR fifo\[13\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_139 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold102 fifo\[12\]\[6\] VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 net14 VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__dlygate4sd3_1
X_0608_ fifo\[0\]\[3\] _0223_ VGND VGND VPWR VPWR _0272_ sky130_fd_sc_hd__or2_1
XFILLER_0_13_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold113 fifo\[4\]\[3\] VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__dlygate4sd3_1
Xhold124 fifo\[12\]\[0\] VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__dlygate4sd3_1
X_0539_ fifo\[14\]\[7\] _0205_ _0206_ fifo\[5\]\[7\] VGND VGND VPWR VPWR _0207_ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0890_ _0001_ _0191_ _0189_ _0408_ VGND VGND VPWR VPWR _0439_ sky130_fd_sc_hd__and4_1
XFILLER_0_42_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0873_ _0429_ VGND VGND VPWR VPWR _0430_ sky130_fd_sc_hd__buf_4
XFILLER_0_42_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0942_ net92 net8 _0460_ VGND VGND VPWR VPWR _0468_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_123 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_148 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1072_ clknet_4_10_0_clk _0111_ VGND VGND VPWR VPWR fifo\[9\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0925_ _0458_ VGND VGND VPWR VPWR _0141_ sky130_fd_sc_hd__clkbuf_1
X_0787_ net81 _0324_ _0379_ VGND VGND VPWR VPWR _0382_ sky130_fd_sc_hd__mux2_1
X_0856_ net45 _0315_ _0420_ VGND VGND VPWR VPWR _0421_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold39 fifo\[2\]\[7\] VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__dlygate4sd3_1
Xhold17 fifo\[15\]\[0\] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__dlygate4sd3_1
Xhold28 fifo\[1\]\[5\] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_48 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0710_ _0338_ VGND VGND VPWR VPWR _0046_ sky130_fd_sc_hd__clkbuf_1
X_0641_ fifo\[9\]\[0\] _0208_ _0209_ fifo\[12\]\[0\] VGND VGND VPWR VPWR _0302_ sky130_fd_sc_hd__a22o_1
X_0572_ _0238_ VGND VGND VPWR VPWR _0027_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1055_ clknet_4_3_0_clk _0094_ VGND VGND VPWR VPWR fifo\[7\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_1124_ clknet_4_4_0_clk _0163_ VGND VGND VPWR VPWR fifo\[15\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0908_ _0196_ _0316_ _0192_ _0317_ VGND VGND VPWR VPWR _0449_ sky130_fd_sc_hd__and4b_1
Xoutput18 net18 VGND VGND VPWR VPWR data_out[6] sky130_fd_sc_hd__buf_2
X_0839_ _0411_ VGND VGND VPWR VPWR _0102_ sky130_fd_sc_hd__clkbuf_1
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0624_ _0286_ VGND VGND VPWR VPWR _0023_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_298 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0555_ _0183_ _0176_ _0179_ _0180_ VGND VGND VPWR VPWR _0223_ sky130_fd_sc_hd__or4_4
X_1038_ clknet_4_5_0_clk _0077_ VGND VGND VPWR VPWR fifo\[4\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_1107_ clknet_4_4_0_clk _0146_ VGND VGND VPWR VPWR fifo\[13\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_224 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold103 fifo\[8\]\[6\] VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__dlygate4sd3_1
X_0538_ _0183_ _0179_ tail\[0\] _0173_ VGND VGND VPWR VPWR _0206_ sky130_fd_sc_hd__and4bb_4
Xhold114 fifo\[7\]\[1\] VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold125 fifo\[3\]\[1\] VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__dlygate4sd3_1
X_0607_ fifo\[3\]\[3\] net23 _0219_ fifo\[15\]\[3\] _0270_ VGND VGND VPWR VPWR _0271_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_28_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0941_ _0467_ VGND VGND VPWR VPWR _0148_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0872_ _0196_ _0316_ _0346_ _0408_ VGND VGND VPWR VPWR _0429_ sky130_fd_sc_hd__and4b_1
XFILLER_0_27_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1071_ clknet_4_9_0_clk _0110_ VGND VGND VPWR VPWR fifo\[9\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_0924_ net62 net8 _0450_ VGND VGND VPWR VPWR _0458_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0855_ _0419_ VGND VGND VPWR VPWR _0420_ sky130_fd_sc_hd__clkbuf_4
X_0786_ _0381_ VGND VGND VPWR VPWR _0079_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold29 fifo\[8\]\[0\] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__dlygate4sd3_1
Xhold18 fifo\[9\]\[0\] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_36_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0571_ net18 _0237_ _0172_ VGND VGND VPWR VPWR _0238_ sky130_fd_sc_hd__mux2_1
X_0640_ fifo\[14\]\[0\] _0205_ _0206_ fifo\[5\]\[0\] VGND VGND VPWR VPWR _0301_ sky130_fd_sc_hd__a22o_1
X_1054_ clknet_4_14_0_clk _0093_ VGND VGND VPWR VPWR fifo\[6\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_1123_ clknet_4_6_0_clk _0162_ VGND VGND VPWR VPWR fifo\[15\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_0907_ _0448_ VGND VGND VPWR VPWR _0133_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput19 net19 VGND VGND VPWR VPWR data_out[7] sky130_fd_sc_hd__clkbuf_4
X_0769_ net115 _0324_ _0369_ VGND VGND VPWR VPWR _0372_ sky130_fd_sc_hd__mux2_1
X_0838_ net56 _0315_ _0410_ VGND VGND VPWR VPWR _0411_ sky130_fd_sc_hd__mux2_1
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0554_ fifo\[3\]\[7\] _0217_ _0219_ fifo\[15\]\[7\] _0221_ VGND VGND VPWR VPWR _0222_
+ sky130_fd_sc_hd__a221o_1
X_0623_ net162 _0285_ _0172_ VGND VGND VPWR VPWR _0286_ sky130_fd_sc_hd__mux2_1
X_1106_ clknet_4_1_0_clk _0145_ VGND VGND VPWR VPWR fifo\[13\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1037_ clknet_4_5_0_clk _0076_ VGND VGND VPWR VPWR fifo\[4\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_236 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold104 fifo\[7\]\[3\] VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__dlygate4sd3_1
Xhold126 fifo\[7\]\[2\] VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold115 fifo\[1\]\[0\] VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0537_ tail\[0\] tail\[1\] _0173_ _0183_ VGND VGND VPWR VPWR _0205_ sky130_fd_sc_hd__and4b_4
X_0606_ fifo\[7\]\[3\] _0175_ _0220_ fifo\[10\]\[3\] VGND VGND VPWR VPWR _0270_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0940_ net149 net7 _0460_ VGND VGND VPWR VPWR _0467_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0871_ _0428_ VGND VGND VPWR VPWR _0117_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1070_ clknet_4_14_0_clk _0109_ VGND VGND VPWR VPWR fifo\[8\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0923_ _0457_ VGND VGND VPWR VPWR _0140_ sky130_fd_sc_hd__clkbuf_1
X_0854_ head\[0\] _0190_ _0317_ _0408_ VGND VGND VPWR VPWR _0419_ sky130_fd_sc_hd__and4_1
XFILLER_0_7_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0785_ net82 _0322_ _0379_ VGND VGND VPWR VPWR _0381_ sky130_fd_sc_hd__mux2_1
Xhold19 fifo\[0\]\[3\] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0570_ _0231_ _0233_ _0235_ _0236_ VGND VGND VPWR VPWR _0237_ sky130_fd_sc_hd__o31a_1
X_1122_ clknet_4_0_0_clk _0161_ VGND VGND VPWR VPWR fifo\[15\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_1053_ clknet_4_15_0_clk _0092_ VGND VGND VPWR VPWR fifo\[6\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_0837_ _0409_ VGND VGND VPWR VPWR _0410_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_43_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0906_ net136 net8 _0440_ VGND VGND VPWR VPWR _0448_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0768_ _0371_ VGND VGND VPWR VPWR _0071_ sky130_fd_sc_hd__clkbuf_1
X_0699_ net33 _0330_ _0320_ VGND VGND VPWR VPWR _0331_ sky130_fd_sc_hd__mux2_1
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0553_ fifo\[7\]\[7\] _0175_ _0220_ fifo\[10\]\[7\] VGND VGND VPWR VPWR _0221_ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0622_ _0279_ _0281_ _0283_ _0284_ VGND VGND VPWR VPWR _0285_ sky130_fd_sc_hd__o31a_1
X_1105_ clknet_4_0_0_clk _0144_ VGND VGND VPWR VPWR fifo\[13\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_1036_ clknet_4_4_0_clk _0075_ VGND VGND VPWR VPWR fifo\[4\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold127 tail\[4\] VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__dlygate4sd3_1
Xhold116 fifo\[6\]\[6\] VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__dlygate4sd3_1
Xhold105 fifo\[5\]\[3\] VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0536_ fifo\[1\]\[7\] net25 net24 fifo\[8\]\[7\] VGND VGND VPWR VPWR _0204_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0605_ fifo\[4\]\[3\] _0212_ _0268_ VGND VGND VPWR VPWR _0269_ sky130_fd_sc_hd__a21o_1
XFILLER_0_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1019_ clknet_4_14_0_clk _0058_ VGND VGND VPWR VPWR fifo\[2\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_318 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0519_ head\[3\] head\[2\] VGND VGND VPWR VPWR _0192_ sky130_fd_sc_hd__and2_1
XFILLER_0_39_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0870_ net40 _0334_ _0420_ VGND VGND VPWR VPWR _0428_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_192 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0999_ clknet_4_3_0_clk _0038_ VGND VGND VPWR VPWR fifo\[0\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0922_ net129 net7 _0450_ VGND VGND VPWR VPWR _0457_ sky130_fd_sc_hd__mux2_1
X_0853_ _0418_ VGND VGND VPWR VPWR _0109_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0784_ _0380_ VGND VGND VPWR VPWR _0078_ sky130_fd_sc_hd__clkbuf_1
Xinput1 data_in[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_2
XFILLER_0_36_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_162 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1121_ clknet_4_0_0_clk _0160_ VGND VGND VPWR VPWR fifo\[15\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_1052_ clknet_4_14_0_clk _0091_ VGND VGND VPWR VPWR fifo\[6\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_0836_ _0196_ _0316_ _0317_ _0408_ VGND VGND VPWR VPWR _0409_ sky130_fd_sc_hd__and4b_1
X_0905_ _0447_ VGND VGND VPWR VPWR _0132_ sky130_fd_sc_hd__clkbuf_1
X_0767_ net88 _0322_ _0369_ VGND VGND VPWR VPWR _0371_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0698_ net6 VGND VGND VPWR VPWR _0330_ sky130_fd_sc_hd__clkbuf_4
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0621_ fifo\[0\]\[2\] _0223_ VGND VGND VPWR VPWR _0284_ sky130_fd_sc_hd__or2_1
X_0552_ _0176_ _0180_ _0179_ _0183_ VGND VGND VPWR VPWR _0220_ sky130_fd_sc_hd__and4bb_4
X_1035_ clknet_4_6_0_clk _0074_ VGND VGND VPWR VPWR fifo\[4\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_1104_ clknet_4_1_0_clk _0143_ VGND VGND VPWR VPWR fifo\[13\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_0819_ net50 _0315_ _0399_ VGND VGND VPWR VPWR _0400_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold106 fifo\[10\]\[6\] VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__dlygate4sd3_1
Xhold128 fifo\[10\]\[2\] VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__dlygate4sd3_1
X_0604_ fifo\[11\]\[3\] _0213_ _0214_ fifo\[13\]\[3\] VGND VGND VPWR VPWR _0268_ sky130_fd_sc_hd__a22o_1
Xhold117 fifo\[13\]\[1\] VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0535_ _0176_ tail\[1\] tail\[0\] tail\[3\] VGND VGND VPWR VPWR _0203_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_124 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1018_ clknet_4_8_0_clk _0057_ VGND VGND VPWR VPWR fifo\[2\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_246 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0518_ head\[1\] head\[0\] VGND VGND VPWR VPWR _0191_ sky130_fd_sc_hd__and2_2
XFILLER_0_39_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_70 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0998_ clknet_4_7_0_clk _0037_ _0019_ VGND VGND VPWR VPWR tail\[3\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_33_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0921_ _0456_ VGND VGND VPWR VPWR _0139_ sky130_fd_sc_hd__clkbuf_1
X_0852_ net47 _0334_ _0410_ VGND VGND VPWR VPWR _0418_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_303 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0783_ net87 _0315_ _0379_ VGND VGND VPWR VPWR _0380_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput2 data_in[1] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__buf_2
XFILLER_0_46_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_174 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1051_ clknet_4_14_0_clk _0090_ VGND VGND VPWR VPWR fifo\[6\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_1120_ clknet_4_2_0_clk _0159_ VGND VGND VPWR VPWR fifo\[15\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0904_ net127 net7 _0440_ VGND VGND VPWR VPWR _0447_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0835_ head\[2\] head\[3\] VGND VGND VPWR VPWR _0408_ sky130_fd_sc_hd__and2b_1
XFILLER_0_43_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0766_ _0370_ VGND VGND VPWR VPWR _0070_ sky130_fd_sc_hd__clkbuf_1
X_0697_ _0329_ VGND VGND VPWR VPWR _0042_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0551_ _0218_ VGND VGND VPWR VPWR _0219_ sky130_fd_sc_hd__clkbuf_4
X_0620_ fifo\[3\]\[2\] net23 _0219_ fifo\[15\]\[2\] _0282_ VGND VGND VPWR VPWR _0283_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1034_ clknet_4_1_0_clk _0073_ VGND VGND VPWR VPWR fifo\[4\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_1103_ clknet_4_1_0_clk _0142_ VGND VGND VPWR VPWR fifo\[13\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0818_ _0398_ VGND VGND VPWR VPWR _0399_ sky130_fd_sc_hd__buf_4
X_0749_ _0360_ VGND VGND VPWR VPWR _0063_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold129 head\[4\] VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0534_ tail\[3\] _0173_ tail\[1\] tail\[0\] VGND VGND VPWR VPWR _0202_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_0_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold107 fifo\[3\]\[3\] VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__dlygate4sd3_1
Xhold118 fifo\[15\]\[2\] VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__dlygate4sd3_1
X_0603_ _0263_ _0264_ _0265_ _0266_ VGND VGND VPWR VPWR _0267_ sky130_fd_sc_hd__or4_1
XFILLER_0_48_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1017_ clknet_4_10_0_clk _0056_ VGND VGND VPWR VPWR fifo\[2\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_258 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0517_ _0189_ VGND VGND VPWR VPWR _0190_ sky130_fd_sc_hd__buf_2
XTAP_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0997_ clknet_4_13_0_clk _0036_ _0018_ VGND VGND VPWR VPWR tail\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0920_ net49 net6 _0450_ VGND VGND VPWR VPWR _0456_ sky130_fd_sc_hd__mux2_1
X_0782_ _0378_ VGND VGND VPWR VPWR _0379_ sky130_fd_sc_hd__buf_4
X_0851_ _0417_ VGND VGND VPWR VPWR _0108_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_315 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput3 data_in[2] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__buf_2
XFILLER_0_52_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1050_ clknet_4_8_0_clk _0089_ VGND VGND VPWR VPWR fifo\[6\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_0834_ _0407_ VGND VGND VPWR VPWR _0101_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0903_ _0446_ VGND VGND VPWR VPWR _0131_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0765_ net59 _0315_ _0369_ VGND VGND VPWR VPWR _0370_ sky130_fd_sc_hd__mux2_1
X_0696_ net30 _0328_ _0320_ VGND VGND VPWR VPWR _0329_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0550_ _0183_ _0176_ _0179_ _0180_ VGND VGND VPWR VPWR _0218_ sky130_fd_sc_hd__and4_1
XFILLER_0_33_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1102_ clknet_4_13_0_clk _0141_ VGND VGND VPWR VPWR fifo\[12\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1033_ clknet_4_0_0_clk _0072_ VGND VGND VPWR VPWR fifo\[4\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_0817_ _0001_ _0191_ _0316_ _0367_ VGND VGND VPWR VPWR _0398_ sky130_fd_sc_hd__and4_1
XFILLER_0_33_96 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0679_ _0189_ VGND VGND VPWR VPWR _0316_ sky130_fd_sc_hd__clkbuf_2
X_0748_ net152 _0322_ _0358_ VGND VGND VPWR VPWR _0360_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold108 fifo\[2\]\[2\] VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0533_ fifo\[2\]\[7\] net166 _0199_ fifo\[6\]\[7\] net165 VGND VGND VPWR VPWR _0201_
+ sky130_fd_sc_hd__a221o_1
X_0602_ fifo\[9\]\[3\] _0208_ _0209_ fifo\[12\]\[3\] VGND VGND VPWR VPWR _0266_ sky130_fd_sc_hd__a22o_1
Xhold119 fifo\[10\]\[3\] VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_28_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_148 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1016_ clknet_4_10_0_clk _0055_ VGND VGND VPWR VPWR fifo\[2\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0516_ _0170_ _0188_ net10 VGND VGND VPWR VPWR _0189_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_39_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0996_ clknet_4_13_0_clk _0035_ _0017_ VGND VGND VPWR VPWR tail\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_14_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_140 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0850_ net130 _0332_ _0410_ VGND VGND VPWR VPWR _0417_ sky130_fd_sc_hd__mux2_1
X_0781_ head\[0\] _0190_ _0317_ _0367_ VGND VGND VPWR VPWR _0378_ sky130_fd_sc_hd__and4_1
XFILLER_0_11_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput4 data_in[3] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__buf_2
XFILLER_0_36_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0979_ _0488_ VGND VGND VPWR VPWR _0165_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0833_ net70 _0334_ _0399_ VGND VGND VPWR VPWR _0407_ sky130_fd_sc_hd__mux2_1
X_0902_ net72 net6 _0440_ VGND VGND VPWR VPWR _0446_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0764_ _0368_ VGND VGND VPWR VPWR _0369_ sky130_fd_sc_hd__clkbuf_4
X_0695_ net5 VGND VGND VPWR VPWR _0328_ sky130_fd_sc_hd__buf_2
XFILLER_0_11_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1101_ clknet_4_15_0_clk _0140_ VGND VGND VPWR VPWR fifo\[12\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_1032_ clknet_4_3_0_clk _0071_ VGND VGND VPWR VPWR fifo\[4\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_0816_ _0397_ VGND VGND VPWR VPWR _0093_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0747_ _0359_ VGND VGND VPWR VPWR _0062_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0678_ net1 VGND VGND VPWR VPWR _0315_ sky130_fd_sc_hd__buf_2
Xhold109 fifo\[11\]\[7\] VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__dlygate4sd3_1
X_0601_ fifo\[14\]\[3\] _0205_ _0206_ fifo\[5\]\[3\] VGND VGND VPWR VPWR _0265_ sky130_fd_sc_hd__a22o_1
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0532_ tail\[3\] _0173_ tail\[1\] _0180_ VGND VGND VPWR VPWR _0200_ sky130_fd_sc_hd__nor4_1
XFILLER_0_44_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1015_ clknet_4_11_0_clk _0054_ VGND VGND VPWR VPWR fifo\[2\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0515_ _0171_ VGND VGND VPWR VPWR _0188_ sky130_fd_sc_hd__inv_2
XTAP_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0995_ clknet_4_12_0_clk _0034_ _0016_ VGND VGND VPWR VPWR tail\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_26_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0780_ _0377_ VGND VGND VPWR VPWR _0077_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput5 data_in[4] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__buf_2
XFILLER_0_52_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0978_ net150 net8 _0480_ VGND VGND VPWR VPWR _0488_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0763_ _0196_ _0316_ _0317_ _0367_ VGND VGND VPWR VPWR _0368_ sky130_fd_sc_hd__and4b_1
XFILLER_0_43_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0832_ _0406_ VGND VGND VPWR VPWR _0100_ sky130_fd_sc_hd__clkbuf_1
X_0901_ _0445_ VGND VGND VPWR VPWR _0130_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0694_ _0327_ VGND VGND VPWR VPWR _0041_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap23 _0217_ VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__buf_2
XFILLER_0_25_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_9_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_9_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_48_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1031_ clknet_4_3_0_clk _0070_ VGND VGND VPWR VPWR fifo\[4\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_1100_ clknet_4_9_0_clk _0139_ VGND VGND VPWR VPWR fifo\[12\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0815_ net43 _0334_ _0389_ VGND VGND VPWR VPWR _0397_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0746_ net35 _0315_ _0358_ VGND VGND VPWR VPWR _0359_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0677_ _0313_ VGND VGND VPWR VPWR _0019_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0531_ tail\[3\] tail\[0\] tail\[1\] _0173_ VGND VGND VPWR VPWR _0199_ sky130_fd_sc_hd__and4bb_4
X_0600_ fifo\[1\]\[3\] net164 net163 fifo\[8\]\[3\] VGND VGND VPWR VPWR _0264_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_231 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1014_ clknet_4_14_0_clk _0053_ VGND VGND VPWR VPWR fifo\[1\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_0729_ _0349_ VGND VGND VPWR VPWR _0054_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0514_ _0186_ _0187_ VGND VGND VPWR VPWR _0034_ sky130_fd_sc_hd__nor2_1
XTAP_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0994_ clknet_4_7_0_clk _0033_ _0015_ VGND VGND VPWR VPWR head\[3\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_41_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput6 data_in[5] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__buf_2
XFILLER_0_36_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0977_ _0487_ VGND VGND VPWR VPWR _0164_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0900_ net138 net5 _0440_ VGND VGND VPWR VPWR _0445_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0762_ head\[3\] head\[2\] VGND VGND VPWR VPWR _0367_ sky130_fd_sc_hd__and2b_1
X_0831_ net102 _0332_ _0399_ VGND VGND VPWR VPWR _0406_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0693_ net46 _0326_ _0320_ VGND VGND VPWR VPWR _0327_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1030_ clknet_4_6_0_clk _0069_ VGND VGND VPWR VPWR fifo\[3\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_0814_ _0396_ VGND VGND VPWR VPWR _0092_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0745_ _0357_ VGND VGND VPWR VPWR _0358_ sky130_fd_sc_hd__clkbuf_4
X_0676_ _0313_ VGND VGND VPWR VPWR _0018_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0530_ tail\[3\] _0173_ tail\[0\] tail\[1\] VGND VGND VPWR VPWR _0198_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_21_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_243 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1013_ clknet_4_15_0_clk _0052_ VGND VGND VPWR VPWR fifo\[1\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_0659_ _0313_ VGND VGND VPWR VPWR _0314_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_12_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0728_ net60 _0315_ _0348_ VGND VGND VPWR VPWR _0349_ sky130_fd_sc_hd__mux2_1
Xclkbuf_4_8_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_8_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_7_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_46 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0513_ _0180_ _0172_ VGND VGND VPWR VPWR _0187_ sky130_fd_sc_hd__nor2_1
XTAP_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0993_ clknet_4_13_0_clk _0032_ _0014_ VGND VGND VPWR VPWR head\[2\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput7 data_in[6] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__buf_2
XFILLER_0_52_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0976_ net148 net7 _0480_ VGND VGND VPWR VPWR _0487_ sky130_fd_sc_hd__mux2_1
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0830_ _0405_ VGND VGND VPWR VPWR _0099_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0761_ _0366_ VGND VGND VPWR VPWR _0069_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0692_ net4 VGND VGND VPWR VPWR _0326_ sky130_fd_sc_hd__buf_2
XFILLER_0_19_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0959_ _0477_ VGND VGND VPWR VPWR _0156_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_274 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput10 push VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__buf_1
X_0813_ net143 _0332_ _0389_ VGND VGND VPWR VPWR _0396_ sky130_fd_sc_hd__mux2_1
X_0744_ _0001_ _0191_ _0316_ _0318_ VGND VGND VPWR VPWR _0357_ sky130_fd_sc_hd__and4_1
X_0675_ _0313_ VGND VGND VPWR VPWR _0017_ sky130_fd_sc_hd__inv_2
X_1089_ clknet_4_0_0_clk _0128_ VGND VGND VPWR VPWR fifo\[11\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1012_ clknet_4_11_0_clk _0051_ VGND VGND VPWR VPWR fifo\[1\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0727_ _0347_ VGND VGND VPWR VPWR _0348_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_12_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0658_ net11 VGND VGND VPWR VPWR _0313_ sky130_fd_sc_hd__buf_4
X_0589_ fifo\[9\]\[4\] _0208_ _0209_ fifo\[12\]\[4\] VGND VGND VPWR VPWR _0254_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_58 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0512_ _0179_ _0186_ _0184_ VGND VGND VPWR VPWR _0035_ sky130_fd_sc_hd__o21a_1
XTAP_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0992_ clknet_4_13_0_clk _0031_ _0013_ VGND VGND VPWR VPWR head\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_41_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_4_7_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_7_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_49_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput8 data_in[7] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_52_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0975_ _0486_ VGND VGND VPWR VPWR _0163_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_250 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0760_ net119 _0334_ _0358_ VGND VGND VPWR VPWR _0366_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0691_ _0325_ VGND VGND VPWR VPWR _0040_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0958_ net118 net7 _0470_ VGND VGND VPWR VPWR _0477_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_286 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0889_ _0438_ VGND VGND VPWR VPWR _0125_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0743_ _0356_ VGND VGND VPWR VPWR _0061_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput11 rst VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_24_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0812_ _0395_ VGND VGND VPWR VPWR _0091_ sky130_fd_sc_hd__clkbuf_1
X_0674_ _0313_ VGND VGND VPWR VPWR _0016_ sky130_fd_sc_hd__inv_2
X_1088_ clknet_4_1_0_clk _0127_ VGND VGND VPWR VPWR fifo\[11\]\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1011_ clknet_4_14_0_clk _0050_ VGND VGND VPWR VPWR fifo\[1\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_0726_ _0196_ _0316_ _0318_ _0346_ VGND VGND VPWR VPWR _0347_ sky130_fd_sc_hd__and4b_1
X_0657_ net11 VGND VGND VPWR VPWR _0001_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0588_ fifo\[14\]\[4\] _0205_ _0206_ fifo\[5\]\[4\] VGND VGND VPWR VPWR _0253_ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0511_ _0185_ _0178_ VGND VGND VPWR VPWR _0186_ sky130_fd_sc_hd__nor2_1
XTAP_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0709_ net142 _0315_ _0337_ VGND VGND VPWR VPWR _0338_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0991_ clknet_4_13_0_clk _0030_ _0012_ VGND VGND VPWR VPWR head\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_41_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput9 pop VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0974_ net63 net6 _0480_ VGND VGND VPWR VPWR _0486_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_6_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_6_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_3_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0690_ net42 _0324_ _0320_ VGND VGND VPWR VPWR _0325_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0957_ _0476_ VGND VGND VPWR VPWR _0155_ sky130_fd_sc_hd__clkbuf_1
X_0888_ net114 net8 _0430_ VGND VGND VPWR VPWR _0438_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0673_ _0313_ VGND VGND VPWR VPWR _0015_ sky130_fd_sc_hd__inv_2
X_0742_ net66 _0334_ _0348_ VGND VGND VPWR VPWR _0356_ sky130_fd_sc_hd__mux2_1
X_0811_ net68 _0330_ _0389_ VGND VGND VPWR VPWR _0395_ sky130_fd_sc_hd__mux2_1
X_1087_ clknet_4_1_0_clk _0126_ VGND VGND VPWR VPWR fifo\[11\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1010_ clknet_4_8_0_clk _0049_ VGND VGND VPWR VPWR fifo\[1\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0656_ net9 net20 net22 net10 VGND VGND VPWR VPWR _0000_ sky130_fd_sc_hd__a22o_1
X_0725_ head\[1\] _0001_ VGND VGND VPWR VPWR _0346_ sky130_fd_sc_hd__and2_1
XFILLER_0_8_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0587_ fifo\[1\]\[4\] net164 net163 fifo\[8\]\[4\] VGND VGND VPWR VPWR _0252_ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0510_ _0180_ VGND VGND VPWR VPWR _0185_ sky130_fd_sc_hd__inv_2
XTAP_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1 fifo\[0\]\[0\] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0708_ _0336_ VGND VGND VPWR VPWR _0337_ sky130_fd_sc_hd__clkbuf_4
X_0639_ fifo\[1\]\[0\] net25 net24 fifo\[8\]\[0\] VGND VGND VPWR VPWR _0300_ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_90 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_135 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0990_ clknet_4_7_0_clk _0000_ _0011_ VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_171 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0973_ _0485_ VGND VGND VPWR VPWR _0162_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0956_ net108 net6 _0470_ VGND VGND VPWR VPWR _0476_ sky130_fd_sc_hd__mux2_1
X_0887_ _0437_ VGND VGND VPWR VPWR _0124_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0810_ _0394_ VGND VGND VPWR VPWR _0090_ sky130_fd_sc_hd__clkbuf_1
X_0672_ _0313_ VGND VGND VPWR VPWR _0014_ sky130_fd_sc_hd__inv_2
X_0741_ _0355_ VGND VGND VPWR VPWR _0060_ sky130_fd_sc_hd__clkbuf_1
X_1086_ clknet_4_4_0_clk _0125_ VGND VGND VPWR VPWR fifo\[10\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0939_ _0466_ VGND VGND VPWR VPWR _0147_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_4_5_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_5_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_53_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_119 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0655_ _0312_ VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__buf_1
X_0724_ _0345_ VGND VGND VPWR VPWR _0053_ sky130_fd_sc_hd__clkbuf_1
X_0586_ fifo\[2\]\[4\] net166 _0199_ fifo\[6\]\[4\] net165 VGND VGND VPWR VPWR _0251_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_47_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1069_ clknet_4_15_0_clk _0108_ VGND VGND VPWR VPWR fifo\[8\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2 fifo\[0\]\[6\] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__dlygate4sd3_1
X_0707_ head\[0\] _0190_ _0317_ _0318_ VGND VGND VPWR VPWR _0336_ sky130_fd_sc_hd__and4_1
XFILLER_0_44_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0569_ fifo\[0\]\[6\] _0223_ VGND VGND VPWR VPWR _0236_ sky130_fd_sc_hd__or2_1
X_0638_ fifo\[2\]\[0\] net27 _0199_ fifo\[6\]\[0\] net26 VGND VGND VPWR VPWR _0299_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0972_ net52 net5 _0480_ VGND VGND VPWR VPWR _0485_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0886_ net133 net7 _0430_ VGND VGND VPWR VPWR _0437_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_158 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0955_ _0475_ VGND VGND VPWR VPWR _0154_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_275 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0740_ net78 _0332_ _0348_ VGND VGND VPWR VPWR _0355_ sky130_fd_sc_hd__mux2_1
X_0671_ _0313_ VGND VGND VPWR VPWR _0013_ sky130_fd_sc_hd__inv_2
X_1085_ clknet_4_5_0_clk _0124_ VGND VGND VPWR VPWR fifo\[10\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_0869_ _0427_ VGND VGND VPWR VPWR _0116_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0938_ net93 net6 _0460_ VGND VGND VPWR VPWR _0466_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0723_ net54 _0334_ _0337_ VGND VGND VPWR VPWR _0345_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0654_ _0170_ _0171_ VGND VGND VPWR VPWR _0312_ sky130_fd_sc_hd__and2_1
X_0585_ _0250_ VGND VGND VPWR VPWR _0026_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1068_ clknet_4_11_0_clk _0107_ VGND VGND VPWR VPWR fifo\[8\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3 fifo\[0\]\[4\] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0706_ _0335_ VGND VGND VPWR VPWR _0045_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_4_4_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_4_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_4_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0568_ fifo\[3\]\[6\] _0217_ _0219_ fifo\[15\]\[6\] _0234_ VGND VGND VPWR VPWR _0235_
+ sky130_fd_sc_hd__a221o_1
X_0499_ _0173_ VGND VGND VPWR VPWR _0176_ sky130_fd_sc_hd__buf_2
XFILLER_0_31_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0637_ _0298_ VGND VGND VPWR VPWR _0022_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_82 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0971_ _0484_ VGND VGND VPWR VPWR _0161_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_118 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0885_ _0436_ VGND VGND VPWR VPWR _0123_ sky130_fd_sc_hd__clkbuf_1
X_0954_ net37 net5 _0470_ VGND VGND VPWR VPWR _0475_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_110 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0670_ _0313_ VGND VGND VPWR VPWR _0012_ sky130_fd_sc_hd__inv_2
X_1084_ clknet_4_1_0_clk _0123_ VGND VGND VPWR VPWR fifo\[10\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0799_ _0196_ _0316_ _0346_ _0367_ VGND VGND VPWR VPWR _0388_ sky130_fd_sc_hd__and4b_1
X_0868_ net61 _0332_ _0420_ VGND VGND VPWR VPWR _0427_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0937_ _0465_ VGND VGND VPWR VPWR _0146_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0653_ _0311_ VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_2
X_0722_ _0344_ VGND VGND VPWR VPWR _0052_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0584_ net159 _0249_ _0172_ VGND VGND VPWR VPWR _0250_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1067_ clknet_4_12_0_clk _0106_ VGND VGND VPWR VPWR fifo\[8\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold4 fifo\[0\]\[1\] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0705_ net32 _0334_ _0320_ VGND VGND VPWR VPWR _0335_ sky130_fd_sc_hd__mux2_1
X_0636_ net13 _0297_ _0172_ VGND VGND VPWR VPWR _0298_ sky130_fd_sc_hd__mux2_1
X_0567_ fifo\[7\]\[6\] _0175_ _0220_ fifo\[10\]\[6\] VGND VGND VPWR VPWR _0234_ sky130_fd_sc_hd__a22o_1
X_0498_ _0174_ VGND VGND VPWR VPWR _0175_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_24_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1119_ clknet_4_3_0_clk _0158_ VGND VGND VPWR VPWR fifo\[15\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0619_ fifo\[7\]\[2\] _0175_ _0220_ fifo\[10\]\[2\] VGND VGND VPWR VPWR _0282_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_3_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_3_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0970_ net157 net4 _0480_ VGND VGND VPWR VPWR _0484_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_214 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0953_ _0474_ VGND VGND VPWR VPWR _0153_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0884_ net137 net6 _0430_ VGND VGND VPWR VPWR _0436_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1083_ clknet_4_6_0_clk _0122_ VGND VGND VPWR VPWR fifo\[10\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0936_ net41 net5 _0460_ VGND VGND VPWR VPWR _0465_ sky130_fd_sc_hd__mux2_1
X_0798_ _0387_ VGND VGND VPWR VPWR _0085_ sky130_fd_sc_hd__clkbuf_1
X_0867_ _0426_ VGND VGND VPWR VPWR _0115_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0652_ _0170_ _0188_ VGND VGND VPWR VPWR _0311_ sky130_fd_sc_hd__and2_1
X_0721_ net117 _0332_ _0337_ VGND VGND VPWR VPWR _0344_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0583_ _0243_ _0245_ _0247_ _0248_ VGND VGND VPWR VPWR _0249_ sky130_fd_sc_hd__o31a_1
XFILLER_0_34_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1066_ clknet_4_8_0_clk _0105_ VGND VGND VPWR VPWR fifo\[8\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_0919_ _0455_ VGND VGND VPWR VPWR _0138_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold5 fifo\[0\]\[7\] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0566_ fifo\[4\]\[6\] _0212_ _0232_ VGND VGND VPWR VPWR _0233_ sky130_fd_sc_hd__a21o_1
X_0704_ net8 VGND VGND VPWR VPWR _0334_ sky130_fd_sc_hd__clkbuf_4
X_0635_ _0291_ _0293_ _0295_ _0296_ VGND VGND VPWR VPWR _0297_ sky130_fd_sc_hd__o31a_1
XFILLER_0_20_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0497_ tail\[3\] _0173_ tail\[1\] tail\[0\] VGND VGND VPWR VPWR _0174_ sky130_fd_sc_hd__and4b_1
XFILLER_0_17_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1118_ clknet_4_15_0_clk _0157_ VGND VGND VPWR VPWR fifo\[14\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_1049_ clknet_4_10_0_clk _0088_ VGND VGND VPWR VPWR fifo\[6\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0549_ _0183_ _0176_ _0181_ VGND VGND VPWR VPWR _0217_ sky130_fd_sc_hd__nor3_1
XFILLER_0_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0618_ fifo\[4\]\[2\] _0212_ _0280_ VGND VGND VPWR VPWR _0281_ sky130_fd_sc_hd__a21o_1
XFILLER_0_48_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire3 _0200_ VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0952_ net116 net4 _0470_ VGND VGND VPWR VPWR _0474_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_226 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0883_ _0435_ VGND VGND VPWR VPWR _0122_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_4_2_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_2_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_5_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1082_ clknet_4_0_0_clk _0121_ VGND VGND VPWR VPWR fifo\[10\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0935_ _0464_ VGND VGND VPWR VPWR _0145_ sky130_fd_sc_hd__clkbuf_1
X_0866_ net51 _0330_ _0420_ VGND VGND VPWR VPWR _0426_ sky130_fd_sc_hd__mux2_1
X_0797_ net85 _0334_ _0379_ VGND VGND VPWR VPWR _0387_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_270 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0720_ _0343_ VGND VGND VPWR VPWR _0051_ sky130_fd_sc_hd__clkbuf_1
X_0651_ net154 _0219_ VGND VGND VPWR VPWR _0020_ sky130_fd_sc_hd__xor2_1
X_0582_ fifo\[0\]\[5\] _0223_ VGND VGND VPWR VPWR _0248_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1065_ clknet_4_9_0_clk _0104_ VGND VGND VPWR VPWR fifo\[8\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_310 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0918_ net96 net5 _0450_ VGND VGND VPWR VPWR _0455_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0849_ _0416_ VGND VGND VPWR VPWR _0107_ sky130_fd_sc_hd__clkbuf_1
Xhold6 fifo\[0\]\[5\] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0703_ _0333_ VGND VGND VPWR VPWR _0044_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_310 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0496_ tail\[2\] VGND VGND VPWR VPWR _0173_ sky130_fd_sc_hd__buf_2
X_0565_ fifo\[11\]\[6\] _0213_ _0214_ fifo\[13\]\[6\] VGND VGND VPWR VPWR _0232_ sky130_fd_sc_hd__a22o_1
X_0634_ fifo\[0\]\[1\] _0223_ VGND VGND VPWR VPWR _0296_ sky130_fd_sc_hd__or2_1
XFILLER_0_20_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1117_ clknet_4_15_0_clk _0156_ VGND VGND VPWR VPWR fifo\[14\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1048_ clknet_4_10_0_clk _0087_ VGND VGND VPWR VPWR fifo\[6\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_118 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0548_ fifo\[4\]\[7\] _0212_ _0215_ VGND VGND VPWR VPWR _0216_ sky130_fd_sc_hd__a21o_1
XFILLER_0_0_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0617_ fifo\[11\]\[2\] _0213_ _0214_ fifo\[13\]\[2\] VGND VGND VPWR VPWR _0280_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4 _0198_ VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_224 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0951_ _0473_ VGND VGND VPWR VPWR _0152_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0882_ net53 net5 _0430_ VGND VGND VPWR VPWR _0435_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_84 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1081_ clknet_4_0_0_clk _0120_ VGND VGND VPWR VPWR fifo\[10\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0865_ _0425_ VGND VGND VPWR VPWR _0114_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0934_ net124 net4 _0460_ VGND VGND VPWR VPWR _0464_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0796_ _0386_ VGND VGND VPWR VPWR _0084_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_282 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0650_ _0310_ VGND VGND VPWR VPWR _0021_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0581_ fifo\[3\]\[5\] net23 _0219_ fifo\[15\]\[5\] _0246_ VGND VGND VPWR VPWR _0247_
+ sky130_fd_sc_hd__a221o_1
Xclkbuf_4_1_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_1_0_clk sky130_fd_sc_hd__clkbuf_8
X_1064_ clknet_4_10_0_clk _0103_ VGND VGND VPWR VPWR fifo\[8\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0779_ net105 _0334_ _0369_ VGND VGND VPWR VPWR _0377_ sky130_fd_sc_hd__mux2_1
X_0917_ _0454_ VGND VGND VPWR VPWR _0137_ sky130_fd_sc_hd__clkbuf_1
X_0848_ net73 _0330_ _0410_ VGND VGND VPWR VPWR _0416_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold7 fifo\[3\]\[4\] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0702_ net29 _0332_ _0320_ VGND VGND VPWR VPWR _0333_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0633_ fifo\[3\]\[1\] net23 _0219_ fifo\[15\]\[1\] _0294_ VGND VGND VPWR VPWR _0295_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_20_32 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0495_ _0170_ _0171_ net9 VGND VGND VPWR VPWR _0172_ sky130_fd_sc_hd__a21boi_4
X_0564_ _0227_ _0228_ _0229_ _0230_ VGND VGND VPWR VPWR _0231_ sky130_fd_sc_hd__or4_1
XFILLER_0_45_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1047_ clknet_4_11_0_clk _0086_ VGND VGND VPWR VPWR fifo\[6\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_1116_ clknet_4_11_0_clk _0155_ VGND VGND VPWR VPWR fifo\[14\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_130 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0616_ _0275_ _0276_ _0277_ _0278_ VGND VGND VPWR VPWR _0279_ sky130_fd_sc_hd__or4_1
X_0547_ fifo\[11\]\[7\] _0213_ _0214_ fifo\[13\]\[7\] VGND VGND VPWR VPWR _0215_ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0881_ _0434_ VGND VGND VPWR VPWR _0121_ sky130_fd_sc_hd__clkbuf_1
X_0950_ net101 net3 _0470_ VGND VGND VPWR VPWR _0473_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_96 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1080_ clknet_4_2_0_clk _0119_ VGND VGND VPWR VPWR fifo\[10\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_0795_ net139 _0332_ _0379_ VGND VGND VPWR VPWR _0386_ sky130_fd_sc_hd__mux2_1
X_0864_ net39 _0328_ _0420_ VGND VGND VPWR VPWR _0425_ sky130_fd_sc_hd__mux2_1
X_0933_ _0463_ VGND VGND VPWR VPWR _0144_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_250 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0580_ fifo\[7\]\[5\] _0175_ _0220_ fifo\[10\]\[5\] VGND VGND VPWR VPWR _0246_ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1063_ clknet_4_11_0_clk _0102_ VGND VGND VPWR VPWR fifo\[8\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0916_ net113 net4 _0450_ VGND VGND VPWR VPWR _0454_ sky130_fd_sc_hd__mux2_1
X_0778_ _0376_ VGND VGND VPWR VPWR _0076_ sky130_fd_sc_hd__clkbuf_1
X_0847_ _0415_ VGND VGND VPWR VPWR _0106_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold8 fifo\[3\]\[0\] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__dlygate4sd3_1
X_0701_ net7 VGND VGND VPWR VPWR _0332_ sky130_fd_sc_hd__clkbuf_4
X_0563_ fifo\[9\]\[6\] _0208_ _0209_ fifo\[12\]\[6\] VGND VGND VPWR VPWR _0230_ sky130_fd_sc_hd__a22o_1
X_0632_ fifo\[7\]\[1\] _0175_ _0220_ fifo\[10\]\[1\] VGND VGND VPWR VPWR _0294_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0494_ head\[4\] tail\[4\] VGND VGND VPWR VPWR _0171_ sky130_fd_sc_hd__xnor2_4
X_1046_ clknet_4_15_0_clk _0085_ VGND VGND VPWR VPWR fifo\[5\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1115_ clknet_4_12_0_clk _0154_ VGND VGND VPWR VPWR fifo\[14\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_4_0_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_0_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0546_ _0179_ _0180_ _0183_ _0176_ VGND VGND VPWR VPWR _0214_ sky130_fd_sc_hd__and4b_4
X_0615_ fifo\[9\]\[2\] _0208_ _0209_ fifo\[12\]\[2\] VGND VGND VPWR VPWR _0278_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1029_ clknet_4_5_0_clk _0068_ VGND VGND VPWR VPWR fifo\[3\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0529_ net156 _0193_ VGND VGND VPWR VPWR _0029_ sky130_fd_sc_hd__xor2_1
XTAP_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_64 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0880_ net146 net4 _0430_ VGND VGND VPWR VPWR _0434_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0932_ net126 net3 _0460_ VGND VGND VPWR VPWR _0463_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0863_ _0424_ VGND VGND VPWR VPWR _0113_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0794_ _0385_ VGND VGND VPWR VPWR _0083_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1062_ clknet_4_4_0_clk _0101_ VGND VGND VPWR VPWR fifo\[7\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_99 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0915_ _0453_ VGND VGND VPWR VPWR _0136_ sky130_fd_sc_hd__clkbuf_1
X_0777_ net64 _0332_ _0369_ VGND VGND VPWR VPWR _0376_ sky130_fd_sc_hd__mux2_1
X_0846_ net38 _0328_ _0410_ VGND VGND VPWR VPWR _0415_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold9 fifo\[4\]\[5\] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_37_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0700_ _0331_ VGND VGND VPWR VPWR _0043_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0562_ fifo\[14\]\[6\] _0205_ _0206_ fifo\[5\]\[6\] VGND VGND VPWR VPWR _0229_ sky130_fd_sc_hd__a22o_1
X_0631_ fifo\[4\]\[1\] _0212_ _0292_ VGND VGND VPWR VPWR _0293_ sky130_fd_sc_hd__a21o_1
XFILLER_0_20_56 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0493_ _0166_ _0167_ _0168_ _0169_ VGND VGND VPWR VPWR _0170_ sky130_fd_sc_hd__and4_2
X_1114_ clknet_4_2_0_clk _0153_ VGND VGND VPWR VPWR fifo\[14\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_1045_ clknet_4_15_0_clk _0084_ VGND VGND VPWR VPWR fifo\[5\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0829_ net99 _0330_ _0399_ VGND VGND VPWR VPWR _0405_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0545_ _0176_ _0179_ _0180_ _0183_ VGND VGND VPWR VPWR _0213_ sky130_fd_sc_hd__and4b_4
XFILLER_0_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0614_ fifo\[14\]\[2\] _0205_ _0206_ fifo\[5\]\[2\] VGND VGND VPWR VPWR _0277_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1028_ clknet_4_1_0_clk _0067_ VGND VGND VPWR VPWR fifo\[3\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0528_ _0196_ _0190_ VGND VGND VPWR VPWR _0030_ sky130_fd_sc_hd__xor2_1
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_143 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0862_ net77 _0326_ _0420_ VGND VGND VPWR VPWR _0424_ sky130_fd_sc_hd__mux2_1
X_0931_ _0462_ VGND VGND VPWR VPWR _0143_ sky130_fd_sc_hd__clkbuf_1
X_0793_ net123 _0330_ _0379_ VGND VGND VPWR VPWR _0385_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1061_ clknet_4_5_0_clk _0100_ VGND VGND VPWR VPWR fifo\[7\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0914_ net83 net3 _0450_ VGND VGND VPWR VPWR _0453_ sky130_fd_sc_hd__mux2_1
X_0845_ _0414_ VGND VGND VPWR VPWR _0105_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0776_ _0375_ VGND VGND VPWR VPWR _0075_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_68 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0492_ tail\[0\] head\[0\] VGND VGND VPWR VPWR _0169_ sky130_fd_sc_hd__xnor2_1
X_0561_ fifo\[1\]\[6\] net25 net24 fifo\[8\]\[6\] VGND VGND VPWR VPWR _0228_ sky130_fd_sc_hd__a22o_1
X_0630_ fifo\[11\]\[1\] _0213_ _0214_ fifo\[13\]\[1\] VGND VGND VPWR VPWR _0292_ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1113_ clknet_4_8_0_clk _0152_ VGND VGND VPWR VPWR fifo\[14\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_1044_ clknet_4_11_0_clk _0083_ VGND VGND VPWR VPWR fifo\[5\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_0759_ _0365_ VGND VGND VPWR VPWR _0068_ sky130_fd_sc_hd__clkbuf_1
X_0828_ _0404_ VGND VGND VPWR VPWR _0098_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_144 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0613_ fifo\[1\]\[2\] net164 net163 fifo\[8\]\[2\] VGND VGND VPWR VPWR _0276_ sky130_fd_sc_hd__a22o_1
XFILLER_0_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0544_ _0183_ _0179_ _0185_ _0176_ VGND VGND VPWR VPWR _0212_ sky130_fd_sc_hd__and4bb_4
XFILLER_0_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1027_ clknet_4_6_0_clk _0066_ VGND VGND VPWR VPWR fifo\[3\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold90 fifo\[1\]\[6\] VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0527_ _0191_ _0190_ _0197_ VGND VGND VPWR VPWR _0031_ sky130_fd_sc_hd__a21oi_1
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_272 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0861_ _0423_ VGND VGND VPWR VPWR _0112_ sky130_fd_sc_hd__clkbuf_1
X_0930_ net144 net2 _0460_ VGND VGND VPWR VPWR _0462_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0792_ _0384_ VGND VGND VPWR VPWR _0082_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xwire24 _0203_ VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_49_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1060_ clknet_4_1_0_clk _0099_ VGND VGND VPWR VPWR fifo\[7\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0913_ _0452_ VGND VGND VPWR VPWR _0135_ sky130_fd_sc_hd__clkbuf_1
X_0844_ net95 _0326_ _0410_ VGND VGND VPWR VPWR _0414_ sky130_fd_sc_hd__mux2_1
X_0775_ net36 _0330_ _0369_ VGND VGND VPWR VPWR _0375_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0491_ tail\[1\] head\[1\] VGND VGND VPWR VPWR _0168_ sky130_fd_sc_hd__xnor2_1
X_0560_ fifo\[2\]\[6\] net166 _0199_ fifo\[6\]\[6\] net165 VGND VGND VPWR VPWR _0227_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_45_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1112_ clknet_4_10_0_clk _0151_ VGND VGND VPWR VPWR fifo\[14\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_1043_ clknet_4_12_0_clk _0082_ VGND VGND VPWR VPWR fifo\[5\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0758_ net71 _0332_ _0358_ VGND VGND VPWR VPWR _0365_ sky130_fd_sc_hd__mux2_1
X_0827_ net100 _0328_ _0399_ VGND VGND VPWR VPWR _0404_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0689_ net3 VGND VGND VPWR VPWR _0324_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_34_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0612_ fifo\[2\]\[2\] net27 _0199_ fifo\[6\]\[2\] net26 VGND VGND VPWR VPWR _0275_
+ sky130_fd_sc_hd__a221o_1
X_0543_ _0201_ _0204_ _0207_ _0210_ VGND VGND VPWR VPWR _0211_ sky130_fd_sc_hd__or4_1
XFILLER_0_8_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1026_ clknet_4_0_0_clk _0065_ VGND VGND VPWR VPWR fifo\[3\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold91 fifo\[14\]\[6\] VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__dlygate4sd3_1
Xhold80 fifo\[2\]\[4\] VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0526_ _0196_ _0190_ net160 VGND VGND VPWR VPWR _0197_ sky130_fd_sc_hd__a21oi_1
XTAP_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1009_ clknet_4_8_0_clk _0048_ VGND VGND VPWR VPWR fifo\[1\]\[2\] sky130_fd_sc_hd__dfxtp_1
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_284 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0509_ _0176_ _0184_ VGND VGND VPWR VPWR _0036_ sky130_fd_sc_hd__xnor2_1
XTAP_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0860_ net90 _0324_ _0420_ VGND VGND VPWR VPWR _0423_ sky130_fd_sc_hd__mux2_1
X_0791_ net111 _0328_ _0379_ VGND VGND VPWR VPWR _0384_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire25 _0202_ VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_80 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0989_ clknet_4_7_0_clk _0029_ _0010_ VGND VGND VPWR VPWR head\[4\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_14_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0912_ net58 net2 _0450_ VGND VGND VPWR VPWR _0452_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0843_ _0413_ VGND VGND VPWR VPWR _0104_ sky130_fd_sc_hd__clkbuf_1
X_0774_ _0374_ VGND VGND VPWR VPWR _0074_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_110 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0490_ tail\[3\] head\[3\] VGND VGND VPWR VPWR _0167_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_29_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_cap1 _0203_ VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__dlymetal6s2s_1
X_1042_ clknet_4_2_0_clk _0081_ VGND VGND VPWR VPWR fifo\[5\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_1111_ clknet_4_9_0_clk _0150_ VGND VGND VPWR VPWR fifo\[14\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0826_ _0403_ VGND VGND VPWR VPWR _0097_ sky130_fd_sc_hd__clkbuf_1
X_0688_ _0323_ VGND VGND VPWR VPWR _0039_ sky130_fd_sc_hd__clkbuf_1
X_0757_ _0364_ VGND VGND VPWR VPWR _0067_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_4_15_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_15_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_34_168 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0542_ fifo\[9\]\[7\] _0208_ _0209_ fifo\[12\]\[7\] VGND VGND VPWR VPWR _0210_ sky130_fd_sc_hd__a22o_1
X_0611_ _0274_ VGND VGND VPWR VPWR _0024_ sky130_fd_sc_hd__clkbuf_1
X_1025_ clknet_4_2_0_clk _0064_ VGND VGND VPWR VPWR fifo\[3\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_168 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_91 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0809_ net80 _0328_ _0389_ VGND VGND VPWR VPWR _0394_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold92 fifo\[3\]\[7\] VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__dlygate4sd3_1
Xhold70 fifo\[1\]\[1\] VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__dlygate4sd3_1
Xhold81 fifo\[14\]\[5\] VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_45_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0525_ head\[0\] VGND VGND VPWR VPWR _0196_ sky130_fd_sc_hd__buf_2
XTAP_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1008_ clknet_4_10_0_clk _0047_ VGND VGND VPWR VPWR fifo\[1\]\[1\] sky130_fd_sc_hd__dfxtp_1
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0508_ _0178_ _0181_ VGND VGND VPWR VPWR _0184_ sky130_fd_sc_hd__or2_1
XTAP_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0790_ _0383_ VGND VGND VPWR VPWR _0081_ sky130_fd_sc_hd__clkbuf_1
Xwire26 net165 VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_2
X_0988_ clknet_4_5_0_clk _0028_ _0009_ VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_92 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_314 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0842_ net57 _0324_ _0410_ VGND VGND VPWR VPWR _0413_ sky130_fd_sc_hd__mux2_1
X_0911_ _0451_ VGND VGND VPWR VPWR _0134_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0773_ net48 _0328_ _0369_ VGND VGND VPWR VPWR _0374_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1110_ clknet_4_5_0_clk _0149_ VGND VGND VPWR VPWR fifo\[13\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap2 _0202_ VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__dlymetal6s2s_1
X_1041_ clknet_4_8_0_clk _0080_ VGND VGND VPWR VPWR fifo\[5\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0825_ net131 _0326_ _0399_ VGND VGND VPWR VPWR _0403_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0687_ net31 _0322_ _0320_ VGND VGND VPWR VPWR _0323_ sky130_fd_sc_hd__mux2_1
X_0756_ net98 _0330_ _0358_ VGND VGND VPWR VPWR _0364_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_144 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0541_ _0179_ _0180_ tail\[3\] _0173_ VGND VGND VPWR VPWR _0209_ sky130_fd_sc_hd__and4bb_4
XFILLER_0_0_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0610_ net15 _0273_ _0172_ VGND VGND VPWR VPWR _0274_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1024_ clknet_4_2_0_clk _0063_ VGND VGND VPWR VPWR fifo\[3\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_0808_ _0393_ VGND VGND VPWR VPWR _0089_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0739_ _0354_ VGND VGND VPWR VPWR _0059_ sky130_fd_sc_hd__clkbuf_1
Xhold93 fifo\[3\]\[2\] VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 fifo\[11\]\[0\] VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__dlygate4sd3_1
Xhold60 fifo\[5\]\[0\] VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 fifo\[3\]\[5\] VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_4_14_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_14_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_5_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0524_ _0194_ _0195_ VGND VGND VPWR VPWR _0032_ sky130_fd_sc_hd__nor2_1
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1007_ clknet_4_11_0_clk _0046_ VGND VGND VPWR VPWR fifo\[1\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0507_ _0172_ _0175_ _0182_ _0183_ VGND VGND VPWR VPWR _0037_ sky130_fd_sc_hd__a22o_1
XTAP_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_38 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xwire27 net166 VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_2
X_0987_ clknet_4_6_0_clk _0027_ _0008_ VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_223 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_172 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0841_ _0412_ VGND VGND VPWR VPWR _0103_ sky130_fd_sc_hd__clkbuf_1
X_0772_ _0373_ VGND VGND VPWR VPWR _0073_ sky130_fd_sc_hd__clkbuf_1
X_0910_ net151 net1 _0450_ VGND VGND VPWR VPWR _0451_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1040_ clknet_4_10_0_clk _0079_ VGND VGND VPWR VPWR fifo\[5\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0824_ _0402_ VGND VGND VPWR VPWR _0096_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0755_ _0363_ VGND VGND VPWR VPWR _0066_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0686_ net2 VGND VGND VPWR VPWR _0322_ sky130_fd_sc_hd__buf_2
XFILLER_0_19_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0540_ _0173_ tail\[1\] tail\[0\] tail\[3\] VGND VGND VPWR VPWR _0208_ sky130_fd_sc_hd__and4bb_4
XFILLER_0_0_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1023_ clknet_4_3_0_clk _0062_ VGND VGND VPWR VPWR fifo\[3\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_0807_ net74 _0326_ _0389_ VGND VGND VPWR VPWR _0393_ sky130_fd_sc_hd__mux2_1
X_0738_ net69 _0330_ _0348_ VGND VGND VPWR VPWR _0354_ sky130_fd_sc_hd__mux2_1
X_0669_ _0314_ VGND VGND VPWR VPWR _0011_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold83 fifo\[9\]\[1\] VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__dlygate4sd3_1
Xhold50 fifo\[9\]\[3\] VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__dlygate4sd3_1
Xhold61 fifo\[4\]\[1\] VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 fifo\[11\]\[1\] VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 fifo\[7\]\[5\] VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0523_ _0191_ _0190_ net161 VGND VGND VPWR VPWR _0195_ sky130_fd_sc_hd__a21oi_1
XTAP_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1006_ clknet_4_7_0_clk _0045_ VGND VGND VPWR VPWR fifo\[0\]\[7\] sky130_fd_sc_hd__dfxtp_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0506_ tail\[3\] VGND VGND VPWR VPWR _0183_ sky130_fd_sc_hd__buf_2
XTAP_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_13_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_13_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_55_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0986_ clknet_4_0_0_clk _0026_ _0007_ VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_151 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0771_ net140 _0326_ _0369_ VGND VGND VPWR VPWR _0373_ sky130_fd_sc_hd__mux2_1
X_0840_ net79 _0322_ _0410_ VGND VGND VPWR VPWR _0412_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0969_ _0483_ VGND VGND VPWR VPWR _0160_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0823_ net153 _0324_ _0399_ VGND VGND VPWR VPWR _0402_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0685_ _0321_ VGND VGND VPWR VPWR _0038_ sky130_fd_sc_hd__clkbuf_1
X_0754_ net34 _0328_ _0358_ VGND VGND VPWR VPWR _0363_ sky130_fd_sc_hd__mux2_1
X_1099_ clknet_4_12_0_clk _0138_ VGND VGND VPWR VPWR fifo\[12\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1022_ clknet_4_14_0_clk _0061_ VGND VGND VPWR VPWR fifo\[2\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_0668_ _0314_ VGND VGND VPWR VPWR _0010_ sky130_fd_sc_hd__inv_2
X_0737_ _0353_ VGND VGND VPWR VPWR _0058_ sky130_fd_sc_hd__clkbuf_1
X_0806_ _0392_ VGND VGND VPWR VPWR _0088_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0599_ fifo\[2\]\[3\] net27 _0199_ fifo\[6\]\[3\] net26 VGND VGND VPWR VPWR _0263_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_15_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold40 fifo\[2\]\[3\] VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold51 fifo\[2\]\[6\] VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 fifo\[7\]\[4\] VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 fifo\[1\]\[3\] VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 fifo\[1\]\[2\] VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 fifo\[5\]\[4\] VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0522_ _0190_ _0193_ _0194_ net158 VGND VGND VPWR VPWR _0033_ sky130_fd_sc_hd__o2bb2a_1
XTAP_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1005_ clknet_4_7_0_clk _0044_ VGND VGND VPWR VPWR fifo\[0\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0505_ _0177_ _0178_ _0181_ VGND VGND VPWR VPWR _0182_ sky130_fd_sc_hd__or3_1
XTAP_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

