module fifo (clk,
    empty,
    error,
    full,
    pop,
    push,
    rst,
    data_in,
    data_out);
 input clk;
 output empty;
 output error;
 output full;
 input pop;
 input push;
 input rst;
 input [7:0] data_in;
 output [7:0] data_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire \fifo[0][0] ;
 wire \fifo[0][1] ;
 wire \fifo[0][2] ;
 wire \fifo[0][3] ;
 wire \fifo[0][4] ;
 wire \fifo[0][5] ;
 wire \fifo[0][6] ;
 wire \fifo[0][7] ;
 wire \fifo[10][0] ;
 wire \fifo[10][1] ;
 wire \fifo[10][2] ;
 wire \fifo[10][3] ;
 wire \fifo[10][4] ;
 wire \fifo[10][5] ;
 wire \fifo[10][6] ;
 wire \fifo[10][7] ;
 wire \fifo[11][0] ;
 wire \fifo[11][1] ;
 wire \fifo[11][2] ;
 wire \fifo[11][3] ;
 wire \fifo[11][4] ;
 wire \fifo[11][5] ;
 wire \fifo[11][6] ;
 wire \fifo[11][7] ;
 wire \fifo[12][0] ;
 wire \fifo[12][1] ;
 wire \fifo[12][2] ;
 wire \fifo[12][3] ;
 wire \fifo[12][4] ;
 wire \fifo[12][5] ;
 wire \fifo[12][6] ;
 wire \fifo[12][7] ;
 wire \fifo[13][0] ;
 wire \fifo[13][1] ;
 wire \fifo[13][2] ;
 wire \fifo[13][3] ;
 wire \fifo[13][4] ;
 wire \fifo[13][5] ;
 wire \fifo[13][6] ;
 wire \fifo[13][7] ;
 wire \fifo[14][0] ;
 wire \fifo[14][1] ;
 wire \fifo[14][2] ;
 wire \fifo[14][3] ;
 wire \fifo[14][4] ;
 wire \fifo[14][5] ;
 wire \fifo[14][6] ;
 wire \fifo[14][7] ;
 wire \fifo[15][0] ;
 wire \fifo[15][1] ;
 wire \fifo[15][2] ;
 wire \fifo[15][3] ;
 wire \fifo[15][4] ;
 wire \fifo[15][5] ;
 wire \fifo[15][6] ;
 wire \fifo[15][7] ;
 wire \fifo[1][0] ;
 wire \fifo[1][1] ;
 wire \fifo[1][2] ;
 wire \fifo[1][3] ;
 wire \fifo[1][4] ;
 wire \fifo[1][5] ;
 wire \fifo[1][6] ;
 wire \fifo[1][7] ;
 wire \fifo[2][0] ;
 wire \fifo[2][1] ;
 wire \fifo[2][2] ;
 wire \fifo[2][3] ;
 wire \fifo[2][4] ;
 wire \fifo[2][5] ;
 wire \fifo[2][6] ;
 wire \fifo[2][7] ;
 wire \fifo[3][0] ;
 wire \fifo[3][1] ;
 wire \fifo[3][2] ;
 wire \fifo[3][3] ;
 wire \fifo[3][4] ;
 wire \fifo[3][5] ;
 wire \fifo[3][6] ;
 wire \fifo[3][7] ;
 wire \fifo[4][0] ;
 wire \fifo[4][1] ;
 wire \fifo[4][2] ;
 wire \fifo[4][3] ;
 wire \fifo[4][4] ;
 wire \fifo[4][5] ;
 wire \fifo[4][6] ;
 wire \fifo[4][7] ;
 wire \fifo[5][0] ;
 wire \fifo[5][1] ;
 wire \fifo[5][2] ;
 wire \fifo[5][3] ;
 wire \fifo[5][4] ;
 wire \fifo[5][5] ;
 wire \fifo[5][6] ;
 wire \fifo[5][7] ;
 wire \fifo[6][0] ;
 wire \fifo[6][1] ;
 wire \fifo[6][2] ;
 wire \fifo[6][3] ;
 wire \fifo[6][4] ;
 wire \fifo[6][5] ;
 wire \fifo[6][6] ;
 wire \fifo[6][7] ;
 wire \fifo[7][0] ;
 wire \fifo[7][1] ;
 wire \fifo[7][2] ;
 wire \fifo[7][3] ;
 wire \fifo[7][4] ;
 wire \fifo[7][5] ;
 wire \fifo[7][6] ;
 wire \fifo[7][7] ;
 wire \fifo[8][0] ;
 wire \fifo[8][1] ;
 wire \fifo[8][2] ;
 wire \fifo[8][3] ;
 wire \fifo[8][4] ;
 wire \fifo[8][5] ;
 wire \fifo[8][6] ;
 wire \fifo[8][7] ;
 wire \fifo[9][0] ;
 wire \fifo[9][1] ;
 wire \fifo[9][2] ;
 wire \fifo[9][3] ;
 wire \fifo[9][4] ;
 wire \fifo[9][5] ;
 wire \fifo[9][6] ;
 wire \fifo[9][7] ;
 wire \head[0] ;
 wire \head[1] ;
 wire \head[2] ;
 wire \head[3] ;
 wire \head[4] ;
 wire \tail[0] ;
 wire \tail[1] ;
 wire \tail[2] ;
 wire \tail[3] ;
 wire \tail[4] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;

 sky130_fd_sc_hd__xnor2_1 _0489_ (.A(\tail[2] ),
    .B(\head[2] ),
    .Y(_0166_));
 sky130_fd_sc_hd__xnor2_1 _0490_ (.A(\tail[3] ),
    .B(\head[3] ),
    .Y(_0167_));
 sky130_fd_sc_hd__xnor2_1 _0491_ (.A(\tail[1] ),
    .B(\head[1] ),
    .Y(_0168_));
 sky130_fd_sc_hd__xnor2_1 _0492_ (.A(\tail[0] ),
    .B(\head[0] ),
    .Y(_0169_));
 sky130_fd_sc_hd__and4_2 _0493_ (.A(_0166_),
    .B(_0167_),
    .C(_0168_),
    .D(_0169_),
    .X(_0170_));
 sky130_fd_sc_hd__xnor2_4 _0494_ (.A(\head[4] ),
    .B(\tail[4] ),
    .Y(_0171_));
 sky130_fd_sc_hd__a21boi_4 _0495_ (.A1(_0170_),
    .A2(_0171_),
    .B1_N(net9),
    .Y(_0172_));
 sky130_fd_sc_hd__buf_2 _0496_ (.A(\tail[2] ),
    .X(_0173_));
 sky130_fd_sc_hd__and4b_1 _0497_ (.A_N(\tail[3] ),
    .B(_0173_),
    .C(\tail[1] ),
    .D(\tail[0] ),
    .X(_0174_));
 sky130_fd_sc_hd__clkbuf_4 _0498_ (.A(_0174_),
    .X(_0175_));
 sky130_fd_sc_hd__buf_2 _0499_ (.A(_0173_),
    .X(_0176_));
 sky130_fd_sc_hd__inv_2 _0500_ (.A(_0176_),
    .Y(_0177_));
 sky130_fd_sc_hd__a21bo_1 _0501_ (.A1(_0170_),
    .A2(_0171_),
    .B1_N(net9),
    .X(_0178_));
 sky130_fd_sc_hd__buf_2 _0502_ (.A(\tail[1] ),
    .X(_0179_));
 sky130_fd_sc_hd__buf_2 _0503_ (.A(\tail[0] ),
    .X(_0180_));
 sky130_fd_sc_hd__nand2_1 _0504_ (.A(_0179_),
    .B(_0180_),
    .Y(_0181_));
 sky130_fd_sc_hd__or3_1 _0505_ (.A(_0177_),
    .B(_0178_),
    .C(_0181_),
    .X(_0182_));
 sky130_fd_sc_hd__buf_2 _0506_ (.A(\tail[3] ),
    .X(_0183_));
 sky130_fd_sc_hd__a22o_1 _0507_ (.A1(_0172_),
    .A2(_0175_),
    .B1(_0182_),
    .B2(_0183_),
    .X(_0037_));
 sky130_fd_sc_hd__or2_1 _0508_ (.A(_0178_),
    .B(_0181_),
    .X(_0184_));
 sky130_fd_sc_hd__xnor2_1 _0509_ (.A(_0176_),
    .B(_0184_),
    .Y(_0036_));
 sky130_fd_sc_hd__inv_2 _0510_ (.A(_0180_),
    .Y(_0185_));
 sky130_fd_sc_hd__nor2_1 _0511_ (.A(_0185_),
    .B(_0178_),
    .Y(_0186_));
 sky130_fd_sc_hd__o21a_1 _0512_ (.A1(_0179_),
    .A2(_0186_),
    .B1(_0184_),
    .X(_0035_));
 sky130_fd_sc_hd__nor2_1 _0513_ (.A(_0180_),
    .B(_0172_),
    .Y(_0187_));
 sky130_fd_sc_hd__nor2_1 _0514_ (.A(_0186_),
    .B(_0187_),
    .Y(_0034_));
 sky130_fd_sc_hd__inv_2 _0515_ (.A(_0171_),
    .Y(_0188_));
 sky130_fd_sc_hd__a21boi_1 _0516_ (.A1(_0170_),
    .A2(_0188_),
    .B1_N(net10),
    .Y(_0189_));
 sky130_fd_sc_hd__buf_2 _0517_ (.A(_0189_),
    .X(_0190_));
 sky130_fd_sc_hd__and2_2 _0518_ (.A(\head[1] ),
    .B(\head[0] ),
    .X(_0191_));
 sky130_fd_sc_hd__and2_1 _0519_ (.A(\head[3] ),
    .B(\head[2] ),
    .X(_0192_));
 sky130_fd_sc_hd__and2_1 _0520_ (.A(_0191_),
    .B(_0192_),
    .X(_0193_));
 sky130_fd_sc_hd__and3_1 _0521_ (.A(\head[2] ),
    .B(_0191_),
    .C(_0190_),
    .X(_0194_));
 sky130_fd_sc_hd__o2bb2a_1 _0522_ (.A1_N(_0190_),
    .A2_N(_0193_),
    .B1(_0194_),
    .B2(net158),
    .X(_0033_));
 sky130_fd_sc_hd__a21oi_1 _0523_ (.A1(_0191_),
    .A2(_0190_),
    .B1(net161),
    .Y(_0195_));
 sky130_fd_sc_hd__nor2_1 _0524_ (.A(_0194_),
    .B(_0195_),
    .Y(_0032_));
 sky130_fd_sc_hd__buf_2 _0525_ (.A(\head[0] ),
    .X(_0196_));
 sky130_fd_sc_hd__a21oi_1 _0526_ (.A1(_0196_),
    .A2(_0190_),
    .B1(net160),
    .Y(_0197_));
 sky130_fd_sc_hd__a21oi_1 _0527_ (.A1(_0191_),
    .A2(_0190_),
    .B1(_0197_),
    .Y(_0031_));
 sky130_fd_sc_hd__xor2_1 _0528_ (.A(_0196_),
    .B(_0190_),
    .X(_0030_));
 sky130_fd_sc_hd__xor2_1 _0529_ (.A(net156),
    .B(_0193_),
    .X(_0029_));
 sky130_fd_sc_hd__nor4b_1 _0530_ (.A(\tail[3] ),
    .B(_0173_),
    .C(\tail[0] ),
    .D_N(\tail[1] ),
    .Y(_0198_));
 sky130_fd_sc_hd__and4bb_4 _0531_ (.A_N(\tail[3] ),
    .B_N(\tail[0] ),
    .C(\tail[1] ),
    .D(_0173_),
    .X(_0199_));
 sky130_fd_sc_hd__nor4_1 _0532_ (.A(\tail[3] ),
    .B(_0173_),
    .C(\tail[1] ),
    .D(_0180_),
    .Y(_0200_));
 sky130_fd_sc_hd__a221o_1 _0533_ (.A1(\fifo[2][7] ),
    .A2(net166),
    .B1(_0199_),
    .B2(\fifo[6][7] ),
    .C1(net165),
    .X(_0201_));
 sky130_fd_sc_hd__nor4b_1 _0534_ (.A(\tail[3] ),
    .B(_0173_),
    .C(\tail[1] ),
    .D_N(\tail[0] ),
    .Y(_0202_));
 sky130_fd_sc_hd__nor4b_1 _0535_ (.A(_0176_),
    .B(\tail[1] ),
    .C(\tail[0] ),
    .D_N(\tail[3] ),
    .Y(_0203_));
 sky130_fd_sc_hd__a22o_1 _0536_ (.A1(\fifo[1][7] ),
    .A2(net25),
    .B1(net24),
    .B2(\fifo[8][7] ),
    .X(_0204_));
 sky130_fd_sc_hd__and4b_4 _0537_ (.A_N(\tail[0] ),
    .B(\tail[1] ),
    .C(_0173_),
    .D(_0183_),
    .X(_0205_));
 sky130_fd_sc_hd__and4bb_4 _0538_ (.A_N(_0183_),
    .B_N(_0179_),
    .C(\tail[0] ),
    .D(_0173_),
    .X(_0206_));
 sky130_fd_sc_hd__a22o_1 _0539_ (.A1(\fifo[14][7] ),
    .A2(_0205_),
    .B1(_0206_),
    .B2(\fifo[5][7] ),
    .X(_0207_));
 sky130_fd_sc_hd__and4bb_4 _0540_ (.A_N(_0173_),
    .B_N(\tail[1] ),
    .C(\tail[0] ),
    .D(\tail[3] ),
    .X(_0208_));
 sky130_fd_sc_hd__and4bb_4 _0541_ (.A_N(_0179_),
    .B_N(_0180_),
    .C(\tail[3] ),
    .D(_0173_),
    .X(_0209_));
 sky130_fd_sc_hd__a22o_1 _0542_ (.A1(\fifo[9][7] ),
    .A2(_0208_),
    .B1(_0209_),
    .B2(\fifo[12][7] ),
    .X(_0210_));
 sky130_fd_sc_hd__or4_1 _0543_ (.A(_0201_),
    .B(_0204_),
    .C(_0207_),
    .D(_0210_),
    .X(_0211_));
 sky130_fd_sc_hd__and4bb_4 _0544_ (.A_N(_0183_),
    .B_N(_0179_),
    .C(_0185_),
    .D(_0176_),
    .X(_0212_));
 sky130_fd_sc_hd__and4b_4 _0545_ (.A_N(_0176_),
    .B(_0179_),
    .C(_0180_),
    .D(_0183_),
    .X(_0213_));
 sky130_fd_sc_hd__and4b_4 _0546_ (.A_N(_0179_),
    .B(_0180_),
    .C(_0183_),
    .D(_0176_),
    .X(_0214_));
 sky130_fd_sc_hd__a22o_1 _0547_ (.A1(\fifo[11][7] ),
    .A2(_0213_),
    .B1(_0214_),
    .B2(\fifo[13][7] ),
    .X(_0215_));
 sky130_fd_sc_hd__a21o_1 _0548_ (.A1(\fifo[4][7] ),
    .A2(_0212_),
    .B1(_0215_),
    .X(_0216_));
 sky130_fd_sc_hd__nor3_1 _0549_ (.A(_0183_),
    .B(_0176_),
    .C(_0181_),
    .Y(_0217_));
 sky130_fd_sc_hd__and4_1 _0550_ (.A(_0183_),
    .B(_0176_),
    .C(_0179_),
    .D(_0180_),
    .X(_0218_));
 sky130_fd_sc_hd__clkbuf_4 _0551_ (.A(_0218_),
    .X(_0219_));
 sky130_fd_sc_hd__and4bb_4 _0552_ (.A_N(_0176_),
    .B_N(_0180_),
    .C(_0179_),
    .D(_0183_),
    .X(_0220_));
 sky130_fd_sc_hd__a22o_1 _0553_ (.A1(\fifo[7][7] ),
    .A2(_0175_),
    .B1(_0220_),
    .B2(\fifo[10][7] ),
    .X(_0221_));
 sky130_fd_sc_hd__a221o_1 _0554_ (.A1(\fifo[3][7] ),
    .A2(_0217_),
    .B1(_0219_),
    .B2(\fifo[15][7] ),
    .C1(_0221_),
    .X(_0222_));
 sky130_fd_sc_hd__or4_4 _0555_ (.A(_0183_),
    .B(_0176_),
    .C(_0179_),
    .D(_0180_),
    .X(_0223_));
 sky130_fd_sc_hd__or2_1 _0556_ (.A(\fifo[0][7] ),
    .B(_0223_),
    .X(_0224_));
 sky130_fd_sc_hd__o31a_1 _0557_ (.A1(_0211_),
    .A2(_0216_),
    .A3(_0222_),
    .B1(_0224_),
    .X(_0225_));
 sky130_fd_sc_hd__mux2_1 _0558_ (.A0(net19),
    .A1(_0225_),
    .S(_0172_),
    .X(_0226_));
 sky130_fd_sc_hd__clkbuf_1 _0559_ (.A(_0226_),
    .X(_0028_));
 sky130_fd_sc_hd__a221o_1 _0560_ (.A1(\fifo[2][6] ),
    .A2(net166),
    .B1(_0199_),
    .B2(\fifo[6][6] ),
    .C1(net165),
    .X(_0227_));
 sky130_fd_sc_hd__a22o_1 _0561_ (.A1(\fifo[1][6] ),
    .A2(net25),
    .B1(net24),
    .B2(\fifo[8][6] ),
    .X(_0228_));
 sky130_fd_sc_hd__a22o_1 _0562_ (.A1(\fifo[14][6] ),
    .A2(_0205_),
    .B1(_0206_),
    .B2(\fifo[5][6] ),
    .X(_0229_));
 sky130_fd_sc_hd__a22o_1 _0563_ (.A1(\fifo[9][6] ),
    .A2(_0208_),
    .B1(_0209_),
    .B2(\fifo[12][6] ),
    .X(_0230_));
 sky130_fd_sc_hd__or4_1 _0564_ (.A(_0227_),
    .B(_0228_),
    .C(_0229_),
    .D(_0230_),
    .X(_0231_));
 sky130_fd_sc_hd__a22o_1 _0565_ (.A1(\fifo[11][6] ),
    .A2(_0213_),
    .B1(_0214_),
    .B2(\fifo[13][6] ),
    .X(_0232_));
 sky130_fd_sc_hd__a21o_1 _0566_ (.A1(\fifo[4][6] ),
    .A2(_0212_),
    .B1(_0232_),
    .X(_0233_));
 sky130_fd_sc_hd__a22o_1 _0567_ (.A1(\fifo[7][6] ),
    .A2(_0175_),
    .B1(_0220_),
    .B2(\fifo[10][6] ),
    .X(_0234_));
 sky130_fd_sc_hd__a221o_1 _0568_ (.A1(\fifo[3][6] ),
    .A2(_0217_),
    .B1(_0219_),
    .B2(\fifo[15][6] ),
    .C1(_0234_),
    .X(_0235_));
 sky130_fd_sc_hd__or2_1 _0569_ (.A(\fifo[0][6] ),
    .B(_0223_),
    .X(_0236_));
 sky130_fd_sc_hd__o31a_1 _0570_ (.A1(_0231_),
    .A2(_0233_),
    .A3(_0235_),
    .B1(_0236_),
    .X(_0237_));
 sky130_fd_sc_hd__mux2_1 _0571_ (.A0(net18),
    .A1(_0237_),
    .S(_0172_),
    .X(_0238_));
 sky130_fd_sc_hd__clkbuf_1 _0572_ (.A(_0238_),
    .X(_0027_));
 sky130_fd_sc_hd__a221o_1 _0573_ (.A1(\fifo[2][5] ),
    .A2(net27),
    .B1(_0199_),
    .B2(\fifo[6][5] ),
    .C1(net26),
    .X(_0239_));
 sky130_fd_sc_hd__a22o_1 _0574_ (.A1(\fifo[1][5] ),
    .A2(net25),
    .B1(net24),
    .B2(\fifo[8][5] ),
    .X(_0240_));
 sky130_fd_sc_hd__a22o_1 _0575_ (.A1(\fifo[14][5] ),
    .A2(_0205_),
    .B1(_0206_),
    .B2(\fifo[5][5] ),
    .X(_0241_));
 sky130_fd_sc_hd__a22o_1 _0576_ (.A1(\fifo[9][5] ),
    .A2(_0208_),
    .B1(_0209_),
    .B2(\fifo[12][5] ),
    .X(_0242_));
 sky130_fd_sc_hd__or4_1 _0577_ (.A(_0239_),
    .B(_0240_),
    .C(_0241_),
    .D(_0242_),
    .X(_0243_));
 sky130_fd_sc_hd__a22o_1 _0578_ (.A1(\fifo[11][5] ),
    .A2(_0213_),
    .B1(_0214_),
    .B2(\fifo[13][5] ),
    .X(_0244_));
 sky130_fd_sc_hd__a21o_1 _0579_ (.A1(\fifo[4][5] ),
    .A2(_0212_),
    .B1(_0244_),
    .X(_0245_));
 sky130_fd_sc_hd__a22o_1 _0580_ (.A1(\fifo[7][5] ),
    .A2(_0175_),
    .B1(_0220_),
    .B2(\fifo[10][5] ),
    .X(_0246_));
 sky130_fd_sc_hd__a221o_1 _0581_ (.A1(\fifo[3][5] ),
    .A2(net23),
    .B1(_0219_),
    .B2(\fifo[15][5] ),
    .C1(_0246_),
    .X(_0247_));
 sky130_fd_sc_hd__or2_1 _0582_ (.A(\fifo[0][5] ),
    .B(_0223_),
    .X(_0248_));
 sky130_fd_sc_hd__o31a_1 _0583_ (.A1(_0243_),
    .A2(_0245_),
    .A3(_0247_),
    .B1(_0248_),
    .X(_0249_));
 sky130_fd_sc_hd__mux2_1 _0584_ (.A0(net159),
    .A1(_0249_),
    .S(_0172_),
    .X(_0250_));
 sky130_fd_sc_hd__clkbuf_1 _0585_ (.A(_0250_),
    .X(_0026_));
 sky130_fd_sc_hd__a221o_1 _0586_ (.A1(\fifo[2][4] ),
    .A2(net166),
    .B1(_0199_),
    .B2(\fifo[6][4] ),
    .C1(net165),
    .X(_0251_));
 sky130_fd_sc_hd__a22o_1 _0587_ (.A1(\fifo[1][4] ),
    .A2(net164),
    .B1(net163),
    .B2(\fifo[8][4] ),
    .X(_0252_));
 sky130_fd_sc_hd__a22o_1 _0588_ (.A1(\fifo[14][4] ),
    .A2(_0205_),
    .B1(_0206_),
    .B2(\fifo[5][4] ),
    .X(_0253_));
 sky130_fd_sc_hd__a22o_1 _0589_ (.A1(\fifo[9][4] ),
    .A2(_0208_),
    .B1(_0209_),
    .B2(\fifo[12][4] ),
    .X(_0254_));
 sky130_fd_sc_hd__or4_1 _0590_ (.A(_0251_),
    .B(_0252_),
    .C(_0253_),
    .D(_0254_),
    .X(_0255_));
 sky130_fd_sc_hd__a22o_1 _0591_ (.A1(\fifo[11][4] ),
    .A2(_0213_),
    .B1(_0214_),
    .B2(\fifo[13][4] ),
    .X(_0256_));
 sky130_fd_sc_hd__a21o_1 _0592_ (.A1(\fifo[4][4] ),
    .A2(_0212_),
    .B1(_0256_),
    .X(_0257_));
 sky130_fd_sc_hd__a22o_1 _0593_ (.A1(\fifo[7][4] ),
    .A2(_0175_),
    .B1(_0220_),
    .B2(\fifo[10][4] ),
    .X(_0258_));
 sky130_fd_sc_hd__a221o_1 _0594_ (.A1(\fifo[3][4] ),
    .A2(net23),
    .B1(_0219_),
    .B2(\fifo[15][4] ),
    .C1(_0258_),
    .X(_0259_));
 sky130_fd_sc_hd__or2_1 _0595_ (.A(\fifo[0][4] ),
    .B(_0223_),
    .X(_0260_));
 sky130_fd_sc_hd__o31a_1 _0596_ (.A1(_0255_),
    .A2(_0257_),
    .A3(_0259_),
    .B1(_0260_),
    .X(_0261_));
 sky130_fd_sc_hd__mux2_1 _0597_ (.A0(net16),
    .A1(_0261_),
    .S(_0172_),
    .X(_0262_));
 sky130_fd_sc_hd__clkbuf_1 _0598_ (.A(_0262_),
    .X(_0025_));
 sky130_fd_sc_hd__a221o_1 _0599_ (.A1(\fifo[2][3] ),
    .A2(net27),
    .B1(_0199_),
    .B2(\fifo[6][3] ),
    .C1(net26),
    .X(_0263_));
 sky130_fd_sc_hd__a22o_1 _0600_ (.A1(\fifo[1][3] ),
    .A2(net164),
    .B1(net163),
    .B2(\fifo[8][3] ),
    .X(_0264_));
 sky130_fd_sc_hd__a22o_1 _0601_ (.A1(\fifo[14][3] ),
    .A2(_0205_),
    .B1(_0206_),
    .B2(\fifo[5][3] ),
    .X(_0265_));
 sky130_fd_sc_hd__a22o_1 _0602_ (.A1(\fifo[9][3] ),
    .A2(_0208_),
    .B1(_0209_),
    .B2(\fifo[12][3] ),
    .X(_0266_));
 sky130_fd_sc_hd__or4_1 _0603_ (.A(_0263_),
    .B(_0264_),
    .C(_0265_),
    .D(_0266_),
    .X(_0267_));
 sky130_fd_sc_hd__a22o_1 _0604_ (.A1(\fifo[11][3] ),
    .A2(_0213_),
    .B1(_0214_),
    .B2(\fifo[13][3] ),
    .X(_0268_));
 sky130_fd_sc_hd__a21o_1 _0605_ (.A1(\fifo[4][3] ),
    .A2(_0212_),
    .B1(_0268_),
    .X(_0269_));
 sky130_fd_sc_hd__a22o_1 _0606_ (.A1(\fifo[7][3] ),
    .A2(_0175_),
    .B1(_0220_),
    .B2(\fifo[10][3] ),
    .X(_0270_));
 sky130_fd_sc_hd__a221o_1 _0607_ (.A1(\fifo[3][3] ),
    .A2(net23),
    .B1(_0219_),
    .B2(\fifo[15][3] ),
    .C1(_0270_),
    .X(_0271_));
 sky130_fd_sc_hd__or2_1 _0608_ (.A(\fifo[0][3] ),
    .B(_0223_),
    .X(_0272_));
 sky130_fd_sc_hd__o31a_1 _0609_ (.A1(_0267_),
    .A2(_0269_),
    .A3(_0271_),
    .B1(_0272_),
    .X(_0273_));
 sky130_fd_sc_hd__mux2_1 _0610_ (.A0(net15),
    .A1(_0273_),
    .S(_0172_),
    .X(_0274_));
 sky130_fd_sc_hd__clkbuf_1 _0611_ (.A(_0274_),
    .X(_0024_));
 sky130_fd_sc_hd__a221o_1 _0612_ (.A1(\fifo[2][2] ),
    .A2(net27),
    .B1(_0199_),
    .B2(\fifo[6][2] ),
    .C1(net26),
    .X(_0275_));
 sky130_fd_sc_hd__a22o_1 _0613_ (.A1(\fifo[1][2] ),
    .A2(net164),
    .B1(net163),
    .B2(\fifo[8][2] ),
    .X(_0276_));
 sky130_fd_sc_hd__a22o_1 _0614_ (.A1(\fifo[14][2] ),
    .A2(_0205_),
    .B1(_0206_),
    .B2(\fifo[5][2] ),
    .X(_0277_));
 sky130_fd_sc_hd__a22o_1 _0615_ (.A1(\fifo[9][2] ),
    .A2(_0208_),
    .B1(_0209_),
    .B2(\fifo[12][2] ),
    .X(_0278_));
 sky130_fd_sc_hd__or4_1 _0616_ (.A(_0275_),
    .B(_0276_),
    .C(_0277_),
    .D(_0278_),
    .X(_0279_));
 sky130_fd_sc_hd__a22o_1 _0617_ (.A1(\fifo[11][2] ),
    .A2(_0213_),
    .B1(_0214_),
    .B2(\fifo[13][2] ),
    .X(_0280_));
 sky130_fd_sc_hd__a21o_1 _0618_ (.A1(\fifo[4][2] ),
    .A2(_0212_),
    .B1(_0280_),
    .X(_0281_));
 sky130_fd_sc_hd__a22o_1 _0619_ (.A1(\fifo[7][2] ),
    .A2(_0175_),
    .B1(_0220_),
    .B2(\fifo[10][2] ),
    .X(_0282_));
 sky130_fd_sc_hd__a221o_1 _0620_ (.A1(\fifo[3][2] ),
    .A2(net23),
    .B1(_0219_),
    .B2(\fifo[15][2] ),
    .C1(_0282_),
    .X(_0283_));
 sky130_fd_sc_hd__or2_1 _0621_ (.A(\fifo[0][2] ),
    .B(_0223_),
    .X(_0284_));
 sky130_fd_sc_hd__o31a_1 _0622_ (.A1(_0279_),
    .A2(_0281_),
    .A3(_0283_),
    .B1(_0284_),
    .X(_0285_));
 sky130_fd_sc_hd__mux2_1 _0623_ (.A0(net162),
    .A1(_0285_),
    .S(_0172_),
    .X(_0286_));
 sky130_fd_sc_hd__clkbuf_1 _0624_ (.A(_0286_),
    .X(_0023_));
 sky130_fd_sc_hd__a221o_1 _0625_ (.A1(\fifo[2][1] ),
    .A2(net27),
    .B1(_0199_),
    .B2(\fifo[6][1] ),
    .C1(net26),
    .X(_0287_));
 sky130_fd_sc_hd__a22o_1 _0626_ (.A1(\fifo[1][1] ),
    .A2(net25),
    .B1(net24),
    .B2(\fifo[8][1] ),
    .X(_0288_));
 sky130_fd_sc_hd__a22o_1 _0627_ (.A1(\fifo[14][1] ),
    .A2(_0205_),
    .B1(_0206_),
    .B2(\fifo[5][1] ),
    .X(_0289_));
 sky130_fd_sc_hd__a22o_1 _0628_ (.A1(\fifo[9][1] ),
    .A2(_0208_),
    .B1(_0209_),
    .B2(\fifo[12][1] ),
    .X(_0290_));
 sky130_fd_sc_hd__or4_1 _0629_ (.A(_0287_),
    .B(_0288_),
    .C(_0289_),
    .D(_0290_),
    .X(_0291_));
 sky130_fd_sc_hd__a22o_1 _0630_ (.A1(\fifo[11][1] ),
    .A2(_0213_),
    .B1(_0214_),
    .B2(\fifo[13][1] ),
    .X(_0292_));
 sky130_fd_sc_hd__a21o_1 _0631_ (.A1(\fifo[4][1] ),
    .A2(_0212_),
    .B1(_0292_),
    .X(_0293_));
 sky130_fd_sc_hd__a22o_1 _0632_ (.A1(\fifo[7][1] ),
    .A2(_0175_),
    .B1(_0220_),
    .B2(\fifo[10][1] ),
    .X(_0294_));
 sky130_fd_sc_hd__a221o_1 _0633_ (.A1(\fifo[3][1] ),
    .A2(net23),
    .B1(_0219_),
    .B2(\fifo[15][1] ),
    .C1(_0294_),
    .X(_0295_));
 sky130_fd_sc_hd__or2_1 _0634_ (.A(\fifo[0][1] ),
    .B(_0223_),
    .X(_0296_));
 sky130_fd_sc_hd__o31a_1 _0635_ (.A1(_0291_),
    .A2(_0293_),
    .A3(_0295_),
    .B1(_0296_),
    .X(_0297_));
 sky130_fd_sc_hd__mux2_1 _0636_ (.A0(net13),
    .A1(_0297_),
    .S(_0172_),
    .X(_0298_));
 sky130_fd_sc_hd__clkbuf_1 _0637_ (.A(_0298_),
    .X(_0022_));
 sky130_fd_sc_hd__a221o_1 _0638_ (.A1(\fifo[2][0] ),
    .A2(net27),
    .B1(_0199_),
    .B2(\fifo[6][0] ),
    .C1(net26),
    .X(_0299_));
 sky130_fd_sc_hd__a22o_1 _0639_ (.A1(\fifo[1][0] ),
    .A2(net25),
    .B1(net24),
    .B2(\fifo[8][0] ),
    .X(_0300_));
 sky130_fd_sc_hd__a22o_1 _0640_ (.A1(\fifo[14][0] ),
    .A2(_0205_),
    .B1(_0206_),
    .B2(\fifo[5][0] ),
    .X(_0301_));
 sky130_fd_sc_hd__a22o_1 _0641_ (.A1(\fifo[9][0] ),
    .A2(_0208_),
    .B1(_0209_),
    .B2(\fifo[12][0] ),
    .X(_0302_));
 sky130_fd_sc_hd__or4_1 _0642_ (.A(_0299_),
    .B(_0300_),
    .C(_0301_),
    .D(_0302_),
    .X(_0303_));
 sky130_fd_sc_hd__a22o_1 _0643_ (.A1(\fifo[11][0] ),
    .A2(_0213_),
    .B1(_0214_),
    .B2(\fifo[13][0] ),
    .X(_0304_));
 sky130_fd_sc_hd__a21o_1 _0644_ (.A1(\fifo[4][0] ),
    .A2(_0212_),
    .B1(_0304_),
    .X(_0305_));
 sky130_fd_sc_hd__a22o_1 _0645_ (.A1(\fifo[7][0] ),
    .A2(_0175_),
    .B1(_0220_),
    .B2(\fifo[10][0] ),
    .X(_0306_));
 sky130_fd_sc_hd__a221o_1 _0646_ (.A1(\fifo[3][0] ),
    .A2(net23),
    .B1(_0219_),
    .B2(\fifo[15][0] ),
    .C1(_0306_),
    .X(_0307_));
 sky130_fd_sc_hd__or2_1 _0647_ (.A(\fifo[0][0] ),
    .B(_0223_),
    .X(_0308_));
 sky130_fd_sc_hd__o31a_1 _0648_ (.A1(_0303_),
    .A2(_0305_),
    .A3(_0307_),
    .B1(_0308_),
    .X(_0309_));
 sky130_fd_sc_hd__mux2_1 _0649_ (.A0(net12),
    .A1(_0309_),
    .S(_0172_),
    .X(_0310_));
 sky130_fd_sc_hd__clkbuf_1 _0650_ (.A(_0310_),
    .X(_0021_));
 sky130_fd_sc_hd__xor2_1 _0651_ (.A(net154),
    .B(_0219_),
    .X(_0020_));
 sky130_fd_sc_hd__and2_1 _0652_ (.A(_0170_),
    .B(_0188_),
    .X(_0311_));
 sky130_fd_sc_hd__clkbuf_2 _0653_ (.A(_0311_),
    .X(net22));
 sky130_fd_sc_hd__and2_1 _0654_ (.A(_0170_),
    .B(_0171_),
    .X(_0312_));
 sky130_fd_sc_hd__buf_1 _0655_ (.A(_0312_),
    .X(net20));
 sky130_fd_sc_hd__a22o_1 _0656_ (.A1(net9),
    .A2(net20),
    .B1(net22),
    .B2(net10),
    .X(_0000_));
 sky130_fd_sc_hd__inv_2 _0657_ (.A(net11),
    .Y(_0001_));
 sky130_fd_sc_hd__buf_4 _0658_ (.A(net11),
    .X(_0313_));
 sky130_fd_sc_hd__clkbuf_8 _0659_ (.A(_0313_),
    .X(_0314_));
 sky130_fd_sc_hd__inv_2 _0660_ (.A(_0314_),
    .Y(_0002_));
 sky130_fd_sc_hd__inv_2 _0661_ (.A(_0314_),
    .Y(_0003_));
 sky130_fd_sc_hd__inv_2 _0662_ (.A(_0314_),
    .Y(_0004_));
 sky130_fd_sc_hd__inv_2 _0663_ (.A(_0314_),
    .Y(_0005_));
 sky130_fd_sc_hd__inv_2 _0664_ (.A(_0314_),
    .Y(_0006_));
 sky130_fd_sc_hd__inv_2 _0665_ (.A(_0314_),
    .Y(_0007_));
 sky130_fd_sc_hd__inv_2 _0666_ (.A(_0314_),
    .Y(_0008_));
 sky130_fd_sc_hd__inv_2 _0667_ (.A(_0314_),
    .Y(_0009_));
 sky130_fd_sc_hd__inv_2 _0668_ (.A(_0314_),
    .Y(_0010_));
 sky130_fd_sc_hd__inv_2 _0669_ (.A(_0314_),
    .Y(_0011_));
 sky130_fd_sc_hd__inv_2 _0670_ (.A(_0313_),
    .Y(_0012_));
 sky130_fd_sc_hd__inv_2 _0671_ (.A(_0313_),
    .Y(_0013_));
 sky130_fd_sc_hd__inv_2 _0672_ (.A(_0313_),
    .Y(_0014_));
 sky130_fd_sc_hd__inv_2 _0673_ (.A(_0313_),
    .Y(_0015_));
 sky130_fd_sc_hd__inv_2 _0674_ (.A(_0313_),
    .Y(_0016_));
 sky130_fd_sc_hd__inv_2 _0675_ (.A(_0313_),
    .Y(_0017_));
 sky130_fd_sc_hd__inv_2 _0676_ (.A(_0313_),
    .Y(_0018_));
 sky130_fd_sc_hd__inv_2 _0677_ (.A(_0313_),
    .Y(_0019_));
 sky130_fd_sc_hd__buf_2 _0678_ (.A(net1),
    .X(_0315_));
 sky130_fd_sc_hd__clkbuf_2 _0679_ (.A(_0189_),
    .X(_0316_));
 sky130_fd_sc_hd__nor2_2 _0680_ (.A(\head[1] ),
    .B(_0313_),
    .Y(_0317_));
 sky130_fd_sc_hd__nor2_1 _0681_ (.A(\head[3] ),
    .B(\head[2] ),
    .Y(_0318_));
 sky130_fd_sc_hd__and4b_1 _0682_ (.A_N(_0196_),
    .B(_0316_),
    .C(_0317_),
    .D(_0318_),
    .X(_0319_));
 sky130_fd_sc_hd__clkbuf_4 _0683_ (.A(_0319_),
    .X(_0320_));
 sky130_fd_sc_hd__mux2_1 _0684_ (.A0(net28),
    .A1(_0315_),
    .S(_0320_),
    .X(_0321_));
 sky130_fd_sc_hd__clkbuf_1 _0685_ (.A(_0321_),
    .X(_0038_));
 sky130_fd_sc_hd__buf_2 _0686_ (.A(net2),
    .X(_0322_));
 sky130_fd_sc_hd__mux2_1 _0687_ (.A0(net31),
    .A1(_0322_),
    .S(_0320_),
    .X(_0323_));
 sky130_fd_sc_hd__clkbuf_1 _0688_ (.A(_0323_),
    .X(_0039_));
 sky130_fd_sc_hd__clkbuf_4 _0689_ (.A(net3),
    .X(_0324_));
 sky130_fd_sc_hd__mux2_1 _0690_ (.A0(net42),
    .A1(_0324_),
    .S(_0320_),
    .X(_0325_));
 sky130_fd_sc_hd__clkbuf_1 _0691_ (.A(_0325_),
    .X(_0040_));
 sky130_fd_sc_hd__buf_2 _0692_ (.A(net4),
    .X(_0326_));
 sky130_fd_sc_hd__mux2_1 _0693_ (.A0(net46),
    .A1(_0326_),
    .S(_0320_),
    .X(_0327_));
 sky130_fd_sc_hd__clkbuf_1 _0694_ (.A(_0327_),
    .X(_0041_));
 sky130_fd_sc_hd__buf_2 _0695_ (.A(net5),
    .X(_0328_));
 sky130_fd_sc_hd__mux2_1 _0696_ (.A0(net30),
    .A1(_0328_),
    .S(_0320_),
    .X(_0329_));
 sky130_fd_sc_hd__clkbuf_1 _0697_ (.A(_0329_),
    .X(_0042_));
 sky130_fd_sc_hd__clkbuf_4 _0698_ (.A(net6),
    .X(_0330_));
 sky130_fd_sc_hd__mux2_1 _0699_ (.A0(net33),
    .A1(_0330_),
    .S(_0320_),
    .X(_0331_));
 sky130_fd_sc_hd__clkbuf_1 _0700_ (.A(_0331_),
    .X(_0043_));
 sky130_fd_sc_hd__clkbuf_4 _0701_ (.A(net7),
    .X(_0332_));
 sky130_fd_sc_hd__mux2_1 _0702_ (.A0(net29),
    .A1(_0332_),
    .S(_0320_),
    .X(_0333_));
 sky130_fd_sc_hd__clkbuf_1 _0703_ (.A(_0333_),
    .X(_0044_));
 sky130_fd_sc_hd__clkbuf_4 _0704_ (.A(net8),
    .X(_0334_));
 sky130_fd_sc_hd__mux2_1 _0705_ (.A0(net32),
    .A1(_0334_),
    .S(_0320_),
    .X(_0335_));
 sky130_fd_sc_hd__clkbuf_1 _0706_ (.A(_0335_),
    .X(_0045_));
 sky130_fd_sc_hd__and4_1 _0707_ (.A(\head[0] ),
    .B(_0190_),
    .C(_0317_),
    .D(_0318_),
    .X(_0336_));
 sky130_fd_sc_hd__clkbuf_4 _0708_ (.A(_0336_),
    .X(_0337_));
 sky130_fd_sc_hd__mux2_1 _0709_ (.A0(net142),
    .A1(_0315_),
    .S(_0337_),
    .X(_0338_));
 sky130_fd_sc_hd__clkbuf_1 _0710_ (.A(_0338_),
    .X(_0046_));
 sky130_fd_sc_hd__mux2_1 _0711_ (.A0(net97),
    .A1(_0322_),
    .S(_0337_),
    .X(_0339_));
 sky130_fd_sc_hd__clkbuf_1 _0712_ (.A(_0339_),
    .X(_0047_));
 sky130_fd_sc_hd__mux2_1 _0713_ (.A0(net89),
    .A1(_0324_),
    .S(_0337_),
    .X(_0340_));
 sky130_fd_sc_hd__clkbuf_1 _0714_ (.A(_0340_),
    .X(_0048_));
 sky130_fd_sc_hd__mux2_1 _0715_ (.A0(net122),
    .A1(_0326_),
    .S(_0337_),
    .X(_0341_));
 sky130_fd_sc_hd__clkbuf_1 _0716_ (.A(_0341_),
    .X(_0049_));
 sky130_fd_sc_hd__mux2_1 _0717_ (.A0(net125),
    .A1(_0328_),
    .S(_0337_),
    .X(_0342_));
 sky130_fd_sc_hd__clkbuf_1 _0718_ (.A(_0342_),
    .X(_0050_));
 sky130_fd_sc_hd__mux2_1 _0719_ (.A0(net55),
    .A1(_0330_),
    .S(_0337_),
    .X(_0343_));
 sky130_fd_sc_hd__clkbuf_1 _0720_ (.A(_0343_),
    .X(_0051_));
 sky130_fd_sc_hd__mux2_1 _0721_ (.A0(net117),
    .A1(_0332_),
    .S(_0337_),
    .X(_0344_));
 sky130_fd_sc_hd__clkbuf_1 _0722_ (.A(_0344_),
    .X(_0052_));
 sky130_fd_sc_hd__mux2_1 _0723_ (.A0(net54),
    .A1(_0334_),
    .S(_0337_),
    .X(_0345_));
 sky130_fd_sc_hd__clkbuf_1 _0724_ (.A(_0345_),
    .X(_0053_));
 sky130_fd_sc_hd__and2_1 _0725_ (.A(\head[1] ),
    .B(_0001_),
    .X(_0346_));
 sky130_fd_sc_hd__and4b_1 _0726_ (.A_N(_0196_),
    .B(_0316_),
    .C(_0318_),
    .D(_0346_),
    .X(_0347_));
 sky130_fd_sc_hd__clkbuf_4 _0727_ (.A(_0347_),
    .X(_0348_));
 sky130_fd_sc_hd__mux2_1 _0728_ (.A0(net60),
    .A1(_0315_),
    .S(_0348_),
    .X(_0349_));
 sky130_fd_sc_hd__clkbuf_1 _0729_ (.A(_0349_),
    .X(_0054_));
 sky130_fd_sc_hd__mux2_1 _0730_ (.A0(net103),
    .A1(_0322_),
    .S(_0348_),
    .X(_0350_));
 sky130_fd_sc_hd__clkbuf_1 _0731_ (.A(_0350_),
    .X(_0055_));
 sky130_fd_sc_hd__mux2_1 _0732_ (.A0(net135),
    .A1(_0324_),
    .S(_0348_),
    .X(_0351_));
 sky130_fd_sc_hd__clkbuf_1 _0733_ (.A(_0351_),
    .X(_0056_));
 sky130_fd_sc_hd__mux2_1 _0734_ (.A0(net67),
    .A1(_0326_),
    .S(_0348_),
    .X(_0352_));
 sky130_fd_sc_hd__clkbuf_1 _0735_ (.A(_0352_),
    .X(_0057_));
 sky130_fd_sc_hd__mux2_1 _0736_ (.A0(net107),
    .A1(_0328_),
    .S(_0348_),
    .X(_0353_));
 sky130_fd_sc_hd__clkbuf_1 _0737_ (.A(_0353_),
    .X(_0058_));
 sky130_fd_sc_hd__mux2_1 _0738_ (.A0(net69),
    .A1(_0330_),
    .S(_0348_),
    .X(_0354_));
 sky130_fd_sc_hd__clkbuf_1 _0739_ (.A(_0354_),
    .X(_0059_));
 sky130_fd_sc_hd__mux2_1 _0740_ (.A0(net78),
    .A1(_0332_),
    .S(_0348_),
    .X(_0355_));
 sky130_fd_sc_hd__clkbuf_1 _0741_ (.A(_0355_),
    .X(_0060_));
 sky130_fd_sc_hd__mux2_1 _0742_ (.A0(net66),
    .A1(_0334_),
    .S(_0348_),
    .X(_0356_));
 sky130_fd_sc_hd__clkbuf_1 _0743_ (.A(_0356_),
    .X(_0061_));
 sky130_fd_sc_hd__and4_1 _0744_ (.A(_0001_),
    .B(_0191_),
    .C(_0316_),
    .D(_0318_),
    .X(_0357_));
 sky130_fd_sc_hd__clkbuf_4 _0745_ (.A(_0357_),
    .X(_0358_));
 sky130_fd_sc_hd__mux2_1 _0746_ (.A0(net35),
    .A1(_0315_),
    .S(_0358_),
    .X(_0359_));
 sky130_fd_sc_hd__clkbuf_1 _0747_ (.A(_0359_),
    .X(_0062_));
 sky130_fd_sc_hd__mux2_1 _0748_ (.A0(net152),
    .A1(_0322_),
    .S(_0358_),
    .X(_0360_));
 sky130_fd_sc_hd__clkbuf_1 _0749_ (.A(_0360_),
    .X(_0063_));
 sky130_fd_sc_hd__mux2_1 _0750_ (.A0(net120),
    .A1(_0324_),
    .S(_0358_),
    .X(_0361_));
 sky130_fd_sc_hd__clkbuf_1 _0751_ (.A(_0361_),
    .X(_0064_));
 sky130_fd_sc_hd__mux2_1 _0752_ (.A0(net134),
    .A1(_0326_),
    .S(_0358_),
    .X(_0362_));
 sky130_fd_sc_hd__clkbuf_1 _0753_ (.A(_0362_),
    .X(_0065_));
 sky130_fd_sc_hd__mux2_1 _0754_ (.A0(net34),
    .A1(_0328_),
    .S(_0358_),
    .X(_0363_));
 sky130_fd_sc_hd__clkbuf_1 _0755_ (.A(_0363_),
    .X(_0066_));
 sky130_fd_sc_hd__mux2_1 _0756_ (.A0(net98),
    .A1(_0330_),
    .S(_0358_),
    .X(_0364_));
 sky130_fd_sc_hd__clkbuf_1 _0757_ (.A(_0364_),
    .X(_0067_));
 sky130_fd_sc_hd__mux2_1 _0758_ (.A0(net71),
    .A1(_0332_),
    .S(_0358_),
    .X(_0365_));
 sky130_fd_sc_hd__clkbuf_1 _0759_ (.A(_0365_),
    .X(_0068_));
 sky130_fd_sc_hd__mux2_1 _0760_ (.A0(net119),
    .A1(_0334_),
    .S(_0358_),
    .X(_0366_));
 sky130_fd_sc_hd__clkbuf_1 _0761_ (.A(_0366_),
    .X(_0069_));
 sky130_fd_sc_hd__and2b_1 _0762_ (.A_N(\head[3] ),
    .B(\head[2] ),
    .X(_0367_));
 sky130_fd_sc_hd__and4b_1 _0763_ (.A_N(_0196_),
    .B(_0316_),
    .C(_0317_),
    .D(_0367_),
    .X(_0368_));
 sky130_fd_sc_hd__clkbuf_4 _0764_ (.A(_0368_),
    .X(_0369_));
 sky130_fd_sc_hd__mux2_1 _0765_ (.A0(net59),
    .A1(_0315_),
    .S(_0369_),
    .X(_0370_));
 sky130_fd_sc_hd__clkbuf_1 _0766_ (.A(_0370_),
    .X(_0070_));
 sky130_fd_sc_hd__mux2_1 _0767_ (.A0(net88),
    .A1(_0322_),
    .S(_0369_),
    .X(_0371_));
 sky130_fd_sc_hd__clkbuf_1 _0768_ (.A(_0371_),
    .X(_0071_));
 sky130_fd_sc_hd__mux2_1 _0769_ (.A0(net115),
    .A1(_0324_),
    .S(_0369_),
    .X(_0372_));
 sky130_fd_sc_hd__clkbuf_1 _0770_ (.A(_0372_),
    .X(_0072_));
 sky130_fd_sc_hd__mux2_1 _0771_ (.A0(net140),
    .A1(_0326_),
    .S(_0369_),
    .X(_0373_));
 sky130_fd_sc_hd__clkbuf_1 _0772_ (.A(_0373_),
    .X(_0073_));
 sky130_fd_sc_hd__mux2_1 _0773_ (.A0(net48),
    .A1(_0328_),
    .S(_0369_),
    .X(_0374_));
 sky130_fd_sc_hd__clkbuf_1 _0774_ (.A(_0374_),
    .X(_0074_));
 sky130_fd_sc_hd__mux2_1 _0775_ (.A0(net36),
    .A1(_0330_),
    .S(_0369_),
    .X(_0375_));
 sky130_fd_sc_hd__clkbuf_1 _0776_ (.A(_0375_),
    .X(_0075_));
 sky130_fd_sc_hd__mux2_1 _0777_ (.A0(net64),
    .A1(_0332_),
    .S(_0369_),
    .X(_0376_));
 sky130_fd_sc_hd__clkbuf_1 _0778_ (.A(_0376_),
    .X(_0076_));
 sky130_fd_sc_hd__mux2_1 _0779_ (.A0(net105),
    .A1(_0334_),
    .S(_0369_),
    .X(_0377_));
 sky130_fd_sc_hd__clkbuf_1 _0780_ (.A(_0377_),
    .X(_0077_));
 sky130_fd_sc_hd__and4_1 _0781_ (.A(\head[0] ),
    .B(_0190_),
    .C(_0317_),
    .D(_0367_),
    .X(_0378_));
 sky130_fd_sc_hd__buf_4 _0782_ (.A(_0378_),
    .X(_0379_));
 sky130_fd_sc_hd__mux2_1 _0783_ (.A0(net87),
    .A1(_0315_),
    .S(_0379_),
    .X(_0380_));
 sky130_fd_sc_hd__clkbuf_1 _0784_ (.A(_0380_),
    .X(_0078_));
 sky130_fd_sc_hd__mux2_1 _0785_ (.A0(net82),
    .A1(_0322_),
    .S(_0379_),
    .X(_0381_));
 sky130_fd_sc_hd__clkbuf_1 _0786_ (.A(_0381_),
    .X(_0079_));
 sky130_fd_sc_hd__mux2_1 _0787_ (.A0(net81),
    .A1(_0324_),
    .S(_0379_),
    .X(_0382_));
 sky130_fd_sc_hd__clkbuf_1 _0788_ (.A(_0382_),
    .X(_0080_));
 sky130_fd_sc_hd__mux2_1 _0789_ (.A0(net132),
    .A1(_0326_),
    .S(_0379_),
    .X(_0383_));
 sky130_fd_sc_hd__clkbuf_1 _0790_ (.A(_0383_),
    .X(_0081_));
 sky130_fd_sc_hd__mux2_1 _0791_ (.A0(net111),
    .A1(_0328_),
    .S(_0379_),
    .X(_0384_));
 sky130_fd_sc_hd__clkbuf_1 _0792_ (.A(_0384_),
    .X(_0082_));
 sky130_fd_sc_hd__mux2_1 _0793_ (.A0(net123),
    .A1(_0330_),
    .S(_0379_),
    .X(_0385_));
 sky130_fd_sc_hd__clkbuf_1 _0794_ (.A(_0385_),
    .X(_0083_));
 sky130_fd_sc_hd__mux2_1 _0795_ (.A0(net139),
    .A1(_0332_),
    .S(_0379_),
    .X(_0386_));
 sky130_fd_sc_hd__clkbuf_1 _0796_ (.A(_0386_),
    .X(_0084_));
 sky130_fd_sc_hd__mux2_1 _0797_ (.A0(net85),
    .A1(_0334_),
    .S(_0379_),
    .X(_0387_));
 sky130_fd_sc_hd__clkbuf_1 _0798_ (.A(_0387_),
    .X(_0085_));
 sky130_fd_sc_hd__and4b_1 _0799_ (.A_N(_0196_),
    .B(_0316_),
    .C(_0346_),
    .D(_0367_),
    .X(_0388_));
 sky130_fd_sc_hd__buf_4 _0800_ (.A(_0388_),
    .X(_0389_));
 sky130_fd_sc_hd__mux2_1 _0801_ (.A0(net75),
    .A1(_0315_),
    .S(_0389_),
    .X(_0390_));
 sky130_fd_sc_hd__clkbuf_1 _0802_ (.A(_0390_),
    .X(_0086_));
 sky130_fd_sc_hd__mux2_1 _0803_ (.A0(net94),
    .A1(_0322_),
    .S(_0389_),
    .X(_0391_));
 sky130_fd_sc_hd__clkbuf_1 _0804_ (.A(_0391_),
    .X(_0087_));
 sky130_fd_sc_hd__mux2_1 _0805_ (.A0(net84),
    .A1(_0324_),
    .S(_0389_),
    .X(_0392_));
 sky130_fd_sc_hd__clkbuf_1 _0806_ (.A(_0392_),
    .X(_0088_));
 sky130_fd_sc_hd__mux2_1 _0807_ (.A0(net74),
    .A1(_0326_),
    .S(_0389_),
    .X(_0393_));
 sky130_fd_sc_hd__clkbuf_1 _0808_ (.A(_0393_),
    .X(_0089_));
 sky130_fd_sc_hd__mux2_1 _0809_ (.A0(net80),
    .A1(_0328_),
    .S(_0389_),
    .X(_0394_));
 sky130_fd_sc_hd__clkbuf_1 _0810_ (.A(_0394_),
    .X(_0090_));
 sky130_fd_sc_hd__mux2_1 _0811_ (.A0(net68),
    .A1(_0330_),
    .S(_0389_),
    .X(_0395_));
 sky130_fd_sc_hd__clkbuf_1 _0812_ (.A(_0395_),
    .X(_0091_));
 sky130_fd_sc_hd__mux2_1 _0813_ (.A0(net143),
    .A1(_0332_),
    .S(_0389_),
    .X(_0396_));
 sky130_fd_sc_hd__clkbuf_1 _0814_ (.A(_0396_),
    .X(_0092_));
 sky130_fd_sc_hd__mux2_1 _0815_ (.A0(net43),
    .A1(_0334_),
    .S(_0389_),
    .X(_0397_));
 sky130_fd_sc_hd__clkbuf_1 _0816_ (.A(_0397_),
    .X(_0093_));
 sky130_fd_sc_hd__and4_1 _0817_ (.A(_0001_),
    .B(_0191_),
    .C(_0316_),
    .D(_0367_),
    .X(_0398_));
 sky130_fd_sc_hd__buf_4 _0818_ (.A(_0398_),
    .X(_0399_));
 sky130_fd_sc_hd__mux2_1 _0819_ (.A0(net50),
    .A1(_0315_),
    .S(_0399_),
    .X(_0400_));
 sky130_fd_sc_hd__clkbuf_1 _0820_ (.A(_0400_),
    .X(_0094_));
 sky130_fd_sc_hd__mux2_1 _0821_ (.A0(net141),
    .A1(_0322_),
    .S(_0399_),
    .X(_0401_));
 sky130_fd_sc_hd__clkbuf_1 _0822_ (.A(_0401_),
    .X(_0095_));
 sky130_fd_sc_hd__mux2_1 _0823_ (.A0(net153),
    .A1(_0324_),
    .S(_0399_),
    .X(_0402_));
 sky130_fd_sc_hd__clkbuf_1 _0824_ (.A(_0402_),
    .X(_0096_));
 sky130_fd_sc_hd__mux2_1 _0825_ (.A0(net131),
    .A1(_0326_),
    .S(_0399_),
    .X(_0403_));
 sky130_fd_sc_hd__clkbuf_1 _0826_ (.A(_0403_),
    .X(_0097_));
 sky130_fd_sc_hd__mux2_1 _0827_ (.A0(net100),
    .A1(_0328_),
    .S(_0399_),
    .X(_0404_));
 sky130_fd_sc_hd__clkbuf_1 _0828_ (.A(_0404_),
    .X(_0098_));
 sky130_fd_sc_hd__mux2_1 _0829_ (.A0(net99),
    .A1(_0330_),
    .S(_0399_),
    .X(_0405_));
 sky130_fd_sc_hd__clkbuf_1 _0830_ (.A(_0405_),
    .X(_0099_));
 sky130_fd_sc_hd__mux2_1 _0831_ (.A0(net102),
    .A1(_0332_),
    .S(_0399_),
    .X(_0406_));
 sky130_fd_sc_hd__clkbuf_1 _0832_ (.A(_0406_),
    .X(_0100_));
 sky130_fd_sc_hd__mux2_1 _0833_ (.A0(net70),
    .A1(_0334_),
    .S(_0399_),
    .X(_0407_));
 sky130_fd_sc_hd__clkbuf_1 _0834_ (.A(_0407_),
    .X(_0101_));
 sky130_fd_sc_hd__and2b_1 _0835_ (.A_N(\head[2] ),
    .B(\head[3] ),
    .X(_0408_));
 sky130_fd_sc_hd__and4b_1 _0836_ (.A_N(_0196_),
    .B(_0316_),
    .C(_0317_),
    .D(_0408_),
    .X(_0409_));
 sky130_fd_sc_hd__clkbuf_4 _0837_ (.A(_0409_),
    .X(_0410_));
 sky130_fd_sc_hd__mux2_1 _0838_ (.A0(net56),
    .A1(_0315_),
    .S(_0410_),
    .X(_0411_));
 sky130_fd_sc_hd__clkbuf_1 _0839_ (.A(_0411_),
    .X(_0102_));
 sky130_fd_sc_hd__mux2_1 _0840_ (.A0(net79),
    .A1(_0322_),
    .S(_0410_),
    .X(_0412_));
 sky130_fd_sc_hd__clkbuf_1 _0841_ (.A(_0412_),
    .X(_0103_));
 sky130_fd_sc_hd__mux2_1 _0842_ (.A0(net57),
    .A1(_0324_),
    .S(_0410_),
    .X(_0413_));
 sky130_fd_sc_hd__clkbuf_1 _0843_ (.A(_0413_),
    .X(_0104_));
 sky130_fd_sc_hd__mux2_1 _0844_ (.A0(net95),
    .A1(_0326_),
    .S(_0410_),
    .X(_0414_));
 sky130_fd_sc_hd__clkbuf_1 _0845_ (.A(_0414_),
    .X(_0105_));
 sky130_fd_sc_hd__mux2_1 _0846_ (.A0(net38),
    .A1(_0328_),
    .S(_0410_),
    .X(_0415_));
 sky130_fd_sc_hd__clkbuf_1 _0847_ (.A(_0415_),
    .X(_0106_));
 sky130_fd_sc_hd__mux2_1 _0848_ (.A0(net73),
    .A1(_0330_),
    .S(_0410_),
    .X(_0416_));
 sky130_fd_sc_hd__clkbuf_1 _0849_ (.A(_0416_),
    .X(_0107_));
 sky130_fd_sc_hd__mux2_1 _0850_ (.A0(net130),
    .A1(_0332_),
    .S(_0410_),
    .X(_0417_));
 sky130_fd_sc_hd__clkbuf_1 _0851_ (.A(_0417_),
    .X(_0108_));
 sky130_fd_sc_hd__mux2_1 _0852_ (.A0(net47),
    .A1(_0334_),
    .S(_0410_),
    .X(_0418_));
 sky130_fd_sc_hd__clkbuf_1 _0853_ (.A(_0418_),
    .X(_0109_));
 sky130_fd_sc_hd__and4_1 _0854_ (.A(\head[0] ),
    .B(_0190_),
    .C(_0317_),
    .D(_0408_),
    .X(_0419_));
 sky130_fd_sc_hd__clkbuf_4 _0855_ (.A(_0419_),
    .X(_0420_));
 sky130_fd_sc_hd__mux2_1 _0856_ (.A0(net45),
    .A1(_0315_),
    .S(_0420_),
    .X(_0421_));
 sky130_fd_sc_hd__clkbuf_1 _0857_ (.A(_0421_),
    .X(_0110_));
 sky130_fd_sc_hd__mux2_1 _0858_ (.A0(net110),
    .A1(_0322_),
    .S(_0420_),
    .X(_0422_));
 sky130_fd_sc_hd__clkbuf_1 _0859_ (.A(_0422_),
    .X(_0111_));
 sky130_fd_sc_hd__mux2_1 _0860_ (.A0(net90),
    .A1(_0324_),
    .S(_0420_),
    .X(_0423_));
 sky130_fd_sc_hd__clkbuf_1 _0861_ (.A(_0423_),
    .X(_0112_));
 sky130_fd_sc_hd__mux2_1 _0862_ (.A0(net77),
    .A1(_0326_),
    .S(_0420_),
    .X(_0424_));
 sky130_fd_sc_hd__clkbuf_1 _0863_ (.A(_0424_),
    .X(_0113_));
 sky130_fd_sc_hd__mux2_1 _0864_ (.A0(net39),
    .A1(_0328_),
    .S(_0420_),
    .X(_0425_));
 sky130_fd_sc_hd__clkbuf_1 _0865_ (.A(_0425_),
    .X(_0114_));
 sky130_fd_sc_hd__mux2_1 _0866_ (.A0(net51),
    .A1(_0330_),
    .S(_0420_),
    .X(_0426_));
 sky130_fd_sc_hd__clkbuf_1 _0867_ (.A(_0426_),
    .X(_0115_));
 sky130_fd_sc_hd__mux2_1 _0868_ (.A0(net61),
    .A1(_0332_),
    .S(_0420_),
    .X(_0427_));
 sky130_fd_sc_hd__clkbuf_1 _0869_ (.A(_0427_),
    .X(_0116_));
 sky130_fd_sc_hd__mux2_1 _0870_ (.A0(net40),
    .A1(_0334_),
    .S(_0420_),
    .X(_0428_));
 sky130_fd_sc_hd__clkbuf_1 _0871_ (.A(_0428_),
    .X(_0117_));
 sky130_fd_sc_hd__and4b_1 _0872_ (.A_N(_0196_),
    .B(_0316_),
    .C(_0346_),
    .D(_0408_),
    .X(_0429_));
 sky130_fd_sc_hd__buf_4 _0873_ (.A(_0429_),
    .X(_0430_));
 sky130_fd_sc_hd__mux2_1 _0874_ (.A0(net104),
    .A1(net1),
    .S(_0430_),
    .X(_0431_));
 sky130_fd_sc_hd__clkbuf_1 _0875_ (.A(_0431_),
    .X(_0118_));
 sky130_fd_sc_hd__mux2_1 _0876_ (.A0(net76),
    .A1(net2),
    .S(_0430_),
    .X(_0432_));
 sky130_fd_sc_hd__clkbuf_1 _0877_ (.A(_0432_),
    .X(_0119_));
 sky130_fd_sc_hd__mux2_1 _0878_ (.A0(net155),
    .A1(net3),
    .S(_0430_),
    .X(_0433_));
 sky130_fd_sc_hd__clkbuf_1 _0879_ (.A(_0433_),
    .X(_0120_));
 sky130_fd_sc_hd__mux2_1 _0880_ (.A0(net146),
    .A1(net4),
    .S(_0430_),
    .X(_0434_));
 sky130_fd_sc_hd__clkbuf_1 _0881_ (.A(_0434_),
    .X(_0121_));
 sky130_fd_sc_hd__mux2_1 _0882_ (.A0(net53),
    .A1(net5),
    .S(_0430_),
    .X(_0435_));
 sky130_fd_sc_hd__clkbuf_1 _0883_ (.A(_0435_),
    .X(_0122_));
 sky130_fd_sc_hd__mux2_1 _0884_ (.A0(net137),
    .A1(net6),
    .S(_0430_),
    .X(_0436_));
 sky130_fd_sc_hd__clkbuf_1 _0885_ (.A(_0436_),
    .X(_0123_));
 sky130_fd_sc_hd__mux2_1 _0886_ (.A0(net133),
    .A1(net7),
    .S(_0430_),
    .X(_0437_));
 sky130_fd_sc_hd__clkbuf_1 _0887_ (.A(_0437_),
    .X(_0124_));
 sky130_fd_sc_hd__mux2_1 _0888_ (.A0(net114),
    .A1(net8),
    .S(_0430_),
    .X(_0438_));
 sky130_fd_sc_hd__clkbuf_1 _0889_ (.A(_0438_),
    .X(_0125_));
 sky130_fd_sc_hd__and4_1 _0890_ (.A(_0001_),
    .B(_0191_),
    .C(_0189_),
    .D(_0408_),
    .X(_0439_));
 sky130_fd_sc_hd__clkbuf_4 _0891_ (.A(_0439_),
    .X(_0440_));
 sky130_fd_sc_hd__mux2_1 _0892_ (.A0(net109),
    .A1(net1),
    .S(_0440_),
    .X(_0441_));
 sky130_fd_sc_hd__clkbuf_1 _0893_ (.A(_0441_),
    .X(_0126_));
 sky130_fd_sc_hd__mux2_1 _0894_ (.A0(net121),
    .A1(net2),
    .S(_0440_),
    .X(_0442_));
 sky130_fd_sc_hd__clkbuf_1 _0895_ (.A(_0442_),
    .X(_0127_));
 sky130_fd_sc_hd__mux2_1 _0896_ (.A0(net147),
    .A1(net3),
    .S(_0440_),
    .X(_0443_));
 sky130_fd_sc_hd__clkbuf_1 _0897_ (.A(_0443_),
    .X(_0128_));
 sky130_fd_sc_hd__mux2_1 _0898_ (.A0(net128),
    .A1(net4),
    .S(_0440_),
    .X(_0444_));
 sky130_fd_sc_hd__clkbuf_1 _0899_ (.A(_0444_),
    .X(_0129_));
 sky130_fd_sc_hd__mux2_1 _0900_ (.A0(net138),
    .A1(net5),
    .S(_0440_),
    .X(_0445_));
 sky130_fd_sc_hd__clkbuf_1 _0901_ (.A(_0445_),
    .X(_0130_));
 sky130_fd_sc_hd__mux2_1 _0902_ (.A0(net72),
    .A1(net6),
    .S(_0440_),
    .X(_0446_));
 sky130_fd_sc_hd__clkbuf_1 _0903_ (.A(_0446_),
    .X(_0131_));
 sky130_fd_sc_hd__mux2_1 _0904_ (.A0(net127),
    .A1(net7),
    .S(_0440_),
    .X(_0447_));
 sky130_fd_sc_hd__clkbuf_1 _0905_ (.A(_0447_),
    .X(_0132_));
 sky130_fd_sc_hd__mux2_1 _0906_ (.A0(net136),
    .A1(net8),
    .S(_0440_),
    .X(_0448_));
 sky130_fd_sc_hd__clkbuf_1 _0907_ (.A(_0448_),
    .X(_0133_));
 sky130_fd_sc_hd__and4b_1 _0908_ (.A_N(_0196_),
    .B(_0316_),
    .C(_0192_),
    .D(_0317_),
    .X(_0449_));
 sky130_fd_sc_hd__buf_4 _0909_ (.A(_0449_),
    .X(_0450_));
 sky130_fd_sc_hd__mux2_1 _0910_ (.A0(net151),
    .A1(net1),
    .S(_0450_),
    .X(_0451_));
 sky130_fd_sc_hd__clkbuf_1 _0911_ (.A(_0451_),
    .X(_0134_));
 sky130_fd_sc_hd__mux2_1 _0912_ (.A0(net58),
    .A1(net2),
    .S(_0450_),
    .X(_0452_));
 sky130_fd_sc_hd__clkbuf_1 _0913_ (.A(_0452_),
    .X(_0135_));
 sky130_fd_sc_hd__mux2_1 _0914_ (.A0(net83),
    .A1(net3),
    .S(_0450_),
    .X(_0453_));
 sky130_fd_sc_hd__clkbuf_1 _0915_ (.A(_0453_),
    .X(_0136_));
 sky130_fd_sc_hd__mux2_1 _0916_ (.A0(net113),
    .A1(net4),
    .S(_0450_),
    .X(_0454_));
 sky130_fd_sc_hd__clkbuf_1 _0917_ (.A(_0454_),
    .X(_0137_));
 sky130_fd_sc_hd__mux2_1 _0918_ (.A0(net96),
    .A1(net5),
    .S(_0450_),
    .X(_0455_));
 sky130_fd_sc_hd__clkbuf_1 _0919_ (.A(_0455_),
    .X(_0138_));
 sky130_fd_sc_hd__mux2_1 _0920_ (.A0(net49),
    .A1(net6),
    .S(_0450_),
    .X(_0456_));
 sky130_fd_sc_hd__clkbuf_1 _0921_ (.A(_0456_),
    .X(_0139_));
 sky130_fd_sc_hd__mux2_1 _0922_ (.A0(net129),
    .A1(net7),
    .S(_0450_),
    .X(_0457_));
 sky130_fd_sc_hd__clkbuf_1 _0923_ (.A(_0457_),
    .X(_0140_));
 sky130_fd_sc_hd__mux2_1 _0924_ (.A0(net62),
    .A1(net8),
    .S(_0450_),
    .X(_0458_));
 sky130_fd_sc_hd__clkbuf_1 _0925_ (.A(_0458_),
    .X(_0141_));
 sky130_fd_sc_hd__and4_1 _0926_ (.A(\head[0] ),
    .B(_0190_),
    .C(_0192_),
    .D(_0317_),
    .X(_0459_));
 sky130_fd_sc_hd__clkbuf_4 _0927_ (.A(_0459_),
    .X(_0460_));
 sky130_fd_sc_hd__mux2_1 _0928_ (.A0(net106),
    .A1(net1),
    .S(_0460_),
    .X(_0461_));
 sky130_fd_sc_hd__clkbuf_1 _0929_ (.A(_0461_),
    .X(_0142_));
 sky130_fd_sc_hd__mux2_1 _0930_ (.A0(net144),
    .A1(net2),
    .S(_0460_),
    .X(_0462_));
 sky130_fd_sc_hd__clkbuf_1 _0931_ (.A(_0462_),
    .X(_0143_));
 sky130_fd_sc_hd__mux2_1 _0932_ (.A0(net126),
    .A1(net3),
    .S(_0460_),
    .X(_0463_));
 sky130_fd_sc_hd__clkbuf_1 _0933_ (.A(_0463_),
    .X(_0144_));
 sky130_fd_sc_hd__mux2_1 _0934_ (.A0(net124),
    .A1(net4),
    .S(_0460_),
    .X(_0464_));
 sky130_fd_sc_hd__clkbuf_1 _0935_ (.A(_0464_),
    .X(_0145_));
 sky130_fd_sc_hd__mux2_1 _0936_ (.A0(net41),
    .A1(net5),
    .S(_0460_),
    .X(_0465_));
 sky130_fd_sc_hd__clkbuf_1 _0937_ (.A(_0465_),
    .X(_0146_));
 sky130_fd_sc_hd__mux2_1 _0938_ (.A0(net93),
    .A1(net6),
    .S(_0460_),
    .X(_0466_));
 sky130_fd_sc_hd__clkbuf_1 _0939_ (.A(_0466_),
    .X(_0147_));
 sky130_fd_sc_hd__mux2_1 _0940_ (.A0(net149),
    .A1(net7),
    .S(_0460_),
    .X(_0467_));
 sky130_fd_sc_hd__clkbuf_1 _0941_ (.A(_0467_),
    .X(_0148_));
 sky130_fd_sc_hd__mux2_1 _0942_ (.A0(net92),
    .A1(net8),
    .S(_0460_),
    .X(_0468_));
 sky130_fd_sc_hd__clkbuf_1 _0943_ (.A(_0468_),
    .X(_0149_));
 sky130_fd_sc_hd__and4b_1 _0944_ (.A_N(_0196_),
    .B(_0316_),
    .C(_0192_),
    .D(_0346_),
    .X(_0469_));
 sky130_fd_sc_hd__buf_4 _0945_ (.A(_0469_),
    .X(_0470_));
 sky130_fd_sc_hd__mux2_1 _0946_ (.A0(net65),
    .A1(net1),
    .S(_0470_),
    .X(_0471_));
 sky130_fd_sc_hd__clkbuf_1 _0947_ (.A(_0471_),
    .X(_0150_));
 sky130_fd_sc_hd__mux2_1 _0948_ (.A0(net91),
    .A1(net2),
    .S(_0470_),
    .X(_0472_));
 sky130_fd_sc_hd__clkbuf_1 _0949_ (.A(_0472_),
    .X(_0151_));
 sky130_fd_sc_hd__mux2_1 _0950_ (.A0(net101),
    .A1(net3),
    .S(_0470_),
    .X(_0473_));
 sky130_fd_sc_hd__clkbuf_1 _0951_ (.A(_0473_),
    .X(_0152_));
 sky130_fd_sc_hd__mux2_1 _0952_ (.A0(net116),
    .A1(net4),
    .S(_0470_),
    .X(_0474_));
 sky130_fd_sc_hd__clkbuf_1 _0953_ (.A(_0474_),
    .X(_0153_));
 sky130_fd_sc_hd__mux2_1 _0954_ (.A0(net37),
    .A1(net5),
    .S(_0470_),
    .X(_0475_));
 sky130_fd_sc_hd__clkbuf_1 _0955_ (.A(_0475_),
    .X(_0154_));
 sky130_fd_sc_hd__mux2_1 _0956_ (.A0(net108),
    .A1(net6),
    .S(_0470_),
    .X(_0476_));
 sky130_fd_sc_hd__clkbuf_1 _0957_ (.A(_0476_),
    .X(_0155_));
 sky130_fd_sc_hd__mux2_1 _0958_ (.A0(net118),
    .A1(net7),
    .S(_0470_),
    .X(_0477_));
 sky130_fd_sc_hd__clkbuf_1 _0959_ (.A(_0477_),
    .X(_0156_));
 sky130_fd_sc_hd__mux2_1 _0960_ (.A0(net112),
    .A1(net8),
    .S(_0470_),
    .X(_0478_));
 sky130_fd_sc_hd__clkbuf_1 _0961_ (.A(_0478_),
    .X(_0157_));
 sky130_fd_sc_hd__and4_1 _0962_ (.A(_0001_),
    .B(_0191_),
    .C(_0189_),
    .D(_0192_),
    .X(_0479_));
 sky130_fd_sc_hd__buf_4 _0963_ (.A(_0479_),
    .X(_0480_));
 sky130_fd_sc_hd__mux2_1 _0964_ (.A0(net44),
    .A1(net1),
    .S(_0480_),
    .X(_0481_));
 sky130_fd_sc_hd__clkbuf_1 _0965_ (.A(_0481_),
    .X(_0158_));
 sky130_fd_sc_hd__mux2_1 _0966_ (.A0(net86),
    .A1(net2),
    .S(_0480_),
    .X(_0482_));
 sky130_fd_sc_hd__clkbuf_1 _0967_ (.A(_0482_),
    .X(_0159_));
 sky130_fd_sc_hd__mux2_1 _0968_ (.A0(net145),
    .A1(net3),
    .S(_0480_),
    .X(_0483_));
 sky130_fd_sc_hd__clkbuf_1 _0969_ (.A(_0483_),
    .X(_0160_));
 sky130_fd_sc_hd__mux2_1 _0970_ (.A0(net157),
    .A1(net4),
    .S(_0480_),
    .X(_0484_));
 sky130_fd_sc_hd__clkbuf_1 _0971_ (.A(_0484_),
    .X(_0161_));
 sky130_fd_sc_hd__mux2_1 _0972_ (.A0(net52),
    .A1(net5),
    .S(_0480_),
    .X(_0485_));
 sky130_fd_sc_hd__clkbuf_1 _0973_ (.A(_0485_),
    .X(_0162_));
 sky130_fd_sc_hd__mux2_1 _0974_ (.A0(net63),
    .A1(net6),
    .S(_0480_),
    .X(_0486_));
 sky130_fd_sc_hd__clkbuf_1 _0975_ (.A(_0486_),
    .X(_0163_));
 sky130_fd_sc_hd__mux2_1 _0976_ (.A0(net148),
    .A1(net7),
    .S(_0480_),
    .X(_0487_));
 sky130_fd_sc_hd__clkbuf_1 _0977_ (.A(_0487_),
    .X(_0164_));
 sky130_fd_sc_hd__mux2_1 _0978_ (.A0(net150),
    .A1(net8),
    .S(_0480_),
    .X(_0488_));
 sky130_fd_sc_hd__clkbuf_1 _0979_ (.A(_0488_),
    .X(_0165_));
 sky130_fd_sc_hd__dfrtp_2 _0980_ (.CLK(clknet_4_7_0_clk),
    .D(_0020_),
    .RESET_B(_0001_),
    .Q(\tail[4] ));
 sky130_fd_sc_hd__dfrtp_1 _0981_ (.CLK(clknet_4_2_0_clk),
    .D(_0021_),
    .RESET_B(_0002_),
    .Q(net12));
 sky130_fd_sc_hd__dfrtp_1 _0982_ (.CLK(clknet_4_2_0_clk),
    .D(_0022_),
    .RESET_B(_0003_),
    .Q(net13));
 sky130_fd_sc_hd__dfrtp_1 _0983_ (.CLK(clknet_4_0_0_clk),
    .D(_0023_),
    .RESET_B(_0004_),
    .Q(net14));
 sky130_fd_sc_hd__dfrtp_1 _0984_ (.CLK(clknet_4_1_0_clk),
    .D(_0024_),
    .RESET_B(_0005_),
    .Q(net15));
 sky130_fd_sc_hd__dfrtp_1 _0985_ (.CLK(clknet_4_2_0_clk),
    .D(_0025_),
    .RESET_B(_0006_),
    .Q(net16));
 sky130_fd_sc_hd__dfrtp_1 _0986_ (.CLK(clknet_4_0_0_clk),
    .D(_0026_),
    .RESET_B(_0007_),
    .Q(net17));
 sky130_fd_sc_hd__dfrtp_1 _0987_ (.CLK(clknet_4_6_0_clk),
    .D(_0027_),
    .RESET_B(_0008_),
    .Q(net18));
 sky130_fd_sc_hd__dfrtp_1 _0988_ (.CLK(clknet_4_5_0_clk),
    .D(_0028_),
    .RESET_B(_0009_),
    .Q(net19));
 sky130_fd_sc_hd__dfrtp_2 _0989_ (.CLK(clknet_4_7_0_clk),
    .D(_0029_),
    .RESET_B(_0010_),
    .Q(\head[4] ));
 sky130_fd_sc_hd__dfrtp_1 _0990_ (.CLK(clknet_4_7_0_clk),
    .D(_0000_),
    .RESET_B(_0011_),
    .Q(net21));
 sky130_fd_sc_hd__dfrtp_2 _0991_ (.CLK(clknet_4_13_0_clk),
    .D(_0030_),
    .RESET_B(_0012_),
    .Q(\head[0] ));
 sky130_fd_sc_hd__dfrtp_2 _0992_ (.CLK(clknet_4_13_0_clk),
    .D(_0031_),
    .RESET_B(_0013_),
    .Q(\head[1] ));
 sky130_fd_sc_hd__dfrtp_4 _0993_ (.CLK(clknet_4_13_0_clk),
    .D(_0032_),
    .RESET_B(_0014_),
    .Q(\head[2] ));
 sky130_fd_sc_hd__dfrtp_2 _0994_ (.CLK(clknet_4_7_0_clk),
    .D(_0033_),
    .RESET_B(_0015_),
    .Q(\head[3] ));
 sky130_fd_sc_hd__dfrtp_4 _0995_ (.CLK(clknet_4_12_0_clk),
    .D(_0034_),
    .RESET_B(_0016_),
    .Q(\tail[0] ));
 sky130_fd_sc_hd__dfrtp_4 _0996_ (.CLK(clknet_4_13_0_clk),
    .D(_0035_),
    .RESET_B(_0017_),
    .Q(\tail[1] ));
 sky130_fd_sc_hd__dfrtp_1 _0997_ (.CLK(clknet_4_13_0_clk),
    .D(_0036_),
    .RESET_B(_0018_),
    .Q(\tail[2] ));
 sky130_fd_sc_hd__dfrtp_4 _0998_ (.CLK(clknet_4_7_0_clk),
    .D(_0037_),
    .RESET_B(_0019_),
    .Q(\tail[3] ));
 sky130_fd_sc_hd__dfxtp_1 _0999_ (.CLK(clknet_4_3_0_clk),
    .D(_0038_),
    .Q(\fifo[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1000_ (.CLK(clknet_4_3_0_clk),
    .D(_0039_),
    .Q(\fifo[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1001_ (.CLK(clknet_4_2_0_clk),
    .D(_0040_),
    .Q(\fifo[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1002_ (.CLK(clknet_4_0_0_clk),
    .D(_0041_),
    .Q(\fifo[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1003_ (.CLK(clknet_4_6_0_clk),
    .D(_0042_),
    .Q(\fifo[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1004_ (.CLK(clknet_4_4_0_clk),
    .D(_0043_),
    .Q(\fifo[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1005_ (.CLK(clknet_4_7_0_clk),
    .D(_0044_),
    .Q(\fifo[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1006_ (.CLK(clknet_4_7_0_clk),
    .D(_0045_),
    .Q(\fifo[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1007_ (.CLK(clknet_4_11_0_clk),
    .D(_0046_),
    .Q(\fifo[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1008_ (.CLK(clknet_4_10_0_clk),
    .D(_0047_),
    .Q(\fifo[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1009_ (.CLK(clknet_4_8_0_clk),
    .D(_0048_),
    .Q(\fifo[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1010_ (.CLK(clknet_4_8_0_clk),
    .D(_0049_),
    .Q(\fifo[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1011_ (.CLK(clknet_4_14_0_clk),
    .D(_0050_),
    .Q(\fifo[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1012_ (.CLK(clknet_4_11_0_clk),
    .D(_0051_),
    .Q(\fifo[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1013_ (.CLK(clknet_4_15_0_clk),
    .D(_0052_),
    .Q(\fifo[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1014_ (.CLK(clknet_4_14_0_clk),
    .D(_0053_),
    .Q(\fifo[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1015_ (.CLK(clknet_4_11_0_clk),
    .D(_0054_),
    .Q(\fifo[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1016_ (.CLK(clknet_4_10_0_clk),
    .D(_0055_),
    .Q(\fifo[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1017_ (.CLK(clknet_4_10_0_clk),
    .D(_0056_),
    .Q(\fifo[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1018_ (.CLK(clknet_4_8_0_clk),
    .D(_0057_),
    .Q(\fifo[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1019_ (.CLK(clknet_4_14_0_clk),
    .D(_0058_),
    .Q(\fifo[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1020_ (.CLK(clknet_4_11_0_clk),
    .D(_0059_),
    .Q(\fifo[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1021_ (.CLK(clknet_4_15_0_clk),
    .D(_0060_),
    .Q(\fifo[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1022_ (.CLK(clknet_4_14_0_clk),
    .D(_0061_),
    .Q(\fifo[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1023_ (.CLK(clknet_4_3_0_clk),
    .D(_0062_),
    .Q(\fifo[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1024_ (.CLK(clknet_4_2_0_clk),
    .D(_0063_),
    .Q(\fifo[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1025_ (.CLK(clknet_4_2_0_clk),
    .D(_0064_),
    .Q(\fifo[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1026_ (.CLK(clknet_4_0_0_clk),
    .D(_0065_),
    .Q(\fifo[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1027_ (.CLK(clknet_4_6_0_clk),
    .D(_0066_),
    .Q(\fifo[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1028_ (.CLK(clknet_4_1_0_clk),
    .D(_0067_),
    .Q(\fifo[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1029_ (.CLK(clknet_4_5_0_clk),
    .D(_0068_),
    .Q(\fifo[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1030_ (.CLK(clknet_4_6_0_clk),
    .D(_0069_),
    .Q(\fifo[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1031_ (.CLK(clknet_4_3_0_clk),
    .D(_0070_),
    .Q(\fifo[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1032_ (.CLK(clknet_4_3_0_clk),
    .D(_0071_),
    .Q(\fifo[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1033_ (.CLK(clknet_4_0_0_clk),
    .D(_0072_),
    .Q(\fifo[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1034_ (.CLK(clknet_4_1_0_clk),
    .D(_0073_),
    .Q(\fifo[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1035_ (.CLK(clknet_4_6_0_clk),
    .D(_0074_),
    .Q(\fifo[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1036_ (.CLK(clknet_4_4_0_clk),
    .D(_0075_),
    .Q(\fifo[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1037_ (.CLK(clknet_4_5_0_clk),
    .D(_0076_),
    .Q(\fifo[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1038_ (.CLK(clknet_4_5_0_clk),
    .D(_0077_),
    .Q(\fifo[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1039_ (.CLK(clknet_4_9_0_clk),
    .D(_0078_),
    .Q(\fifo[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1040_ (.CLK(clknet_4_10_0_clk),
    .D(_0079_),
    .Q(\fifo[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1041_ (.CLK(clknet_4_8_0_clk),
    .D(_0080_),
    .Q(\fifo[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1042_ (.CLK(clknet_4_2_0_clk),
    .D(_0081_),
    .Q(\fifo[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1043_ (.CLK(clknet_4_12_0_clk),
    .D(_0082_),
    .Q(\fifo[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1044_ (.CLK(clknet_4_11_0_clk),
    .D(_0083_),
    .Q(\fifo[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1045_ (.CLK(clknet_4_15_0_clk),
    .D(_0084_),
    .Q(\fifo[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1046_ (.CLK(clknet_4_15_0_clk),
    .D(_0085_),
    .Q(\fifo[5][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1047_ (.CLK(clknet_4_11_0_clk),
    .D(_0086_),
    .Q(\fifo[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1048_ (.CLK(clknet_4_10_0_clk),
    .D(_0087_),
    .Q(\fifo[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1049_ (.CLK(clknet_4_10_0_clk),
    .D(_0088_),
    .Q(\fifo[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1050_ (.CLK(clknet_4_8_0_clk),
    .D(_0089_),
    .Q(\fifo[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1051_ (.CLK(clknet_4_14_0_clk),
    .D(_0090_),
    .Q(\fifo[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1052_ (.CLK(clknet_4_14_0_clk),
    .D(_0091_),
    .Q(\fifo[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1053_ (.CLK(clknet_4_15_0_clk),
    .D(_0092_),
    .Q(\fifo[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1054_ (.CLK(clknet_4_14_0_clk),
    .D(_0093_),
    .Q(\fifo[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1055_ (.CLK(clknet_4_3_0_clk),
    .D(_0094_),
    .Q(\fifo[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1056_ (.CLK(clknet_4_2_0_clk),
    .D(_0095_),
    .Q(\fifo[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1057_ (.CLK(clknet_4_0_0_clk),
    .D(_0096_),
    .Q(\fifo[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1058_ (.CLK(clknet_4_0_0_clk),
    .D(_0097_),
    .Q(\fifo[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1059_ (.CLK(clknet_4_6_0_clk),
    .D(_0098_),
    .Q(\fifo[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1060_ (.CLK(clknet_4_1_0_clk),
    .D(_0099_),
    .Q(\fifo[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1061_ (.CLK(clknet_4_5_0_clk),
    .D(_0100_),
    .Q(\fifo[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1062_ (.CLK(clknet_4_4_0_clk),
    .D(_0101_),
    .Q(\fifo[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1063_ (.CLK(clknet_4_11_0_clk),
    .D(_0102_),
    .Q(\fifo[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1064_ (.CLK(clknet_4_10_0_clk),
    .D(_0103_),
    .Q(\fifo[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1065_ (.CLK(clknet_4_9_0_clk),
    .D(_0104_),
    .Q(\fifo[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1066_ (.CLK(clknet_4_8_0_clk),
    .D(_0105_),
    .Q(\fifo[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1067_ (.CLK(clknet_4_12_0_clk),
    .D(_0106_),
    .Q(\fifo[8][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1068_ (.CLK(clknet_4_11_0_clk),
    .D(_0107_),
    .Q(\fifo[8][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1069_ (.CLK(clknet_4_15_0_clk),
    .D(_0108_),
    .Q(\fifo[8][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1070_ (.CLK(clknet_4_14_0_clk),
    .D(_0109_),
    .Q(\fifo[8][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1071_ (.CLK(clknet_4_9_0_clk),
    .D(_0110_),
    .Q(\fifo[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1072_ (.CLK(clknet_4_10_0_clk),
    .D(_0111_),
    .Q(\fifo[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1073_ (.CLK(clknet_4_8_0_clk),
    .D(_0112_),
    .Q(\fifo[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1074_ (.CLK(clknet_4_8_0_clk),
    .D(_0113_),
    .Q(\fifo[9][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1075_ (.CLK(clknet_4_12_0_clk),
    .D(_0114_),
    .Q(\fifo[9][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1076_ (.CLK(clknet_4_9_0_clk),
    .D(_0115_),
    .Q(\fifo[9][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1077_ (.CLK(clknet_4_15_0_clk),
    .D(_0116_),
    .Q(\fifo[9][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1078_ (.CLK(clknet_4_13_0_clk),
    .D(_0117_),
    .Q(\fifo[9][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1079_ (.CLK(clknet_4_1_0_clk),
    .D(_0118_),
    .Q(\fifo[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1080_ (.CLK(clknet_4_2_0_clk),
    .D(_0119_),
    .Q(\fifo[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1081_ (.CLK(clknet_4_0_0_clk),
    .D(_0120_),
    .Q(\fifo[10][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1082_ (.CLK(clknet_4_0_0_clk),
    .D(_0121_),
    .Q(\fifo[10][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1083_ (.CLK(clknet_4_6_0_clk),
    .D(_0122_),
    .Q(\fifo[10][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1084_ (.CLK(clknet_4_1_0_clk),
    .D(_0123_),
    .Q(\fifo[10][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1085_ (.CLK(clknet_4_5_0_clk),
    .D(_0124_),
    .Q(\fifo[10][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1086_ (.CLK(clknet_4_4_0_clk),
    .D(_0125_),
    .Q(\fifo[10][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1087_ (.CLK(clknet_4_1_0_clk),
    .D(_0126_),
    .Q(\fifo[11][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1088_ (.CLK(clknet_4_1_0_clk),
    .D(_0127_),
    .Q(\fifo[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1089_ (.CLK(clknet_4_0_0_clk),
    .D(_0128_),
    .Q(\fifo[11][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1090_ (.CLK(clknet_4_1_0_clk),
    .D(_0129_),
    .Q(\fifo[11][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1091_ (.CLK(clknet_4_4_0_clk),
    .D(_0130_),
    .Q(\fifo[11][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1092_ (.CLK(clknet_4_4_0_clk),
    .D(_0131_),
    .Q(\fifo[11][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1093_ (.CLK(clknet_4_5_0_clk),
    .D(_0132_),
    .Q(\fifo[11][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1094_ (.CLK(clknet_4_5_0_clk),
    .D(_0133_),
    .Q(\fifo[11][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1095_ (.CLK(clknet_4_9_0_clk),
    .D(_0134_),
    .Q(\fifo[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1096_ (.CLK(clknet_4_10_0_clk),
    .D(_0135_),
    .Q(\fifo[12][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1097_ (.CLK(clknet_4_8_0_clk),
    .D(_0136_),
    .Q(\fifo[12][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1098_ (.CLK(clknet_4_2_0_clk),
    .D(_0137_),
    .Q(\fifo[12][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1099_ (.CLK(clknet_4_12_0_clk),
    .D(_0138_),
    .Q(\fifo[12][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1100_ (.CLK(clknet_4_9_0_clk),
    .D(_0139_),
    .Q(\fifo[12][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1101_ (.CLK(clknet_4_15_0_clk),
    .D(_0140_),
    .Q(\fifo[12][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1102_ (.CLK(clknet_4_13_0_clk),
    .D(_0141_),
    .Q(\fifo[12][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1103_ (.CLK(clknet_4_1_0_clk),
    .D(_0142_),
    .Q(\fifo[13][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1104_ (.CLK(clknet_4_1_0_clk),
    .D(_0143_),
    .Q(\fifo[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1105_ (.CLK(clknet_4_0_0_clk),
    .D(_0144_),
    .Q(\fifo[13][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1106_ (.CLK(clknet_4_1_0_clk),
    .D(_0145_),
    .Q(\fifo[13][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1107_ (.CLK(clknet_4_4_0_clk),
    .D(_0146_),
    .Q(\fifo[13][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1108_ (.CLK(clknet_4_4_0_clk),
    .D(_0147_),
    .Q(\fifo[13][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1109_ (.CLK(clknet_4_5_0_clk),
    .D(_0148_),
    .Q(\fifo[13][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1110_ (.CLK(clknet_4_5_0_clk),
    .D(_0149_),
    .Q(\fifo[13][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1111_ (.CLK(clknet_4_9_0_clk),
    .D(_0150_),
    .Q(\fifo[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1112_ (.CLK(clknet_4_10_0_clk),
    .D(_0151_),
    .Q(\fifo[14][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1113_ (.CLK(clknet_4_8_0_clk),
    .D(_0152_),
    .Q(\fifo[14][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1114_ (.CLK(clknet_4_2_0_clk),
    .D(_0153_),
    .Q(\fifo[14][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1115_ (.CLK(clknet_4_12_0_clk),
    .D(_0154_),
    .Q(\fifo[14][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1116_ (.CLK(clknet_4_11_0_clk),
    .D(_0155_),
    .Q(\fifo[14][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1117_ (.CLK(clknet_4_15_0_clk),
    .D(_0156_),
    .Q(\fifo[14][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1118_ (.CLK(clknet_4_15_0_clk),
    .D(_0157_),
    .Q(\fifo[14][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1119_ (.CLK(clknet_4_3_0_clk),
    .D(_0158_),
    .Q(\fifo[15][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1120_ (.CLK(clknet_4_2_0_clk),
    .D(_0159_),
    .Q(\fifo[15][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1121_ (.CLK(clknet_4_0_0_clk),
    .D(_0160_),
    .Q(\fifo[15][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1122_ (.CLK(clknet_4_0_0_clk),
    .D(_0161_),
    .Q(\fifo[15][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1123_ (.CLK(clknet_4_6_0_clk),
    .D(_0162_),
    .Q(\fifo[15][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1124_ (.CLK(clknet_4_4_0_clk),
    .D(_0163_),
    .Q(\fifo[15][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1125_ (.CLK(clknet_4_5_0_clk),
    .D(_0164_),
    .Q(\fifo[15][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1126_ (.CLK(clknet_4_5_0_clk),
    .D(_0165_),
    .Q(\fifo[15][7] ));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__buf_2 input1 (.A(data_in[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_2 input2 (.A(data_in[1]),
    .X(net2));
 sky130_fd_sc_hd__buf_2 input3 (.A(data_in[2]),
    .X(net3));
 sky130_fd_sc_hd__buf_2 input4 (.A(data_in[3]),
    .X(net4));
 sky130_fd_sc_hd__buf_2 input5 (.A(data_in[4]),
    .X(net5));
 sky130_fd_sc_hd__buf_2 input6 (.A(data_in[5]),
    .X(net6));
 sky130_fd_sc_hd__buf_2 input7 (.A(data_in[6]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_4 input8 (.A(data_in[7]),
    .X(net8));
 sky130_fd_sc_hd__dlymetal6s2s_1 input9 (.A(pop),
    .X(net9));
 sky130_fd_sc_hd__buf_1 input10 (.A(push),
    .X(net10));
 sky130_fd_sc_hd__dlymetal6s2s_1 input11 (.A(rst),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_4 output12 (.A(net12),
    .X(data_out[0]));
 sky130_fd_sc_hd__clkbuf_4 output13 (.A(net13),
    .X(data_out[1]));
 sky130_fd_sc_hd__clkbuf_4 output14 (.A(net14),
    .X(data_out[2]));
 sky130_fd_sc_hd__clkbuf_4 output15 (.A(net15),
    .X(data_out[3]));
 sky130_fd_sc_hd__buf_2 output16 (.A(net16),
    .X(data_out[4]));
 sky130_fd_sc_hd__clkbuf_4 output17 (.A(net17),
    .X(data_out[5]));
 sky130_fd_sc_hd__buf_2 output18 (.A(net18),
    .X(data_out[6]));
 sky130_fd_sc_hd__clkbuf_4 output19 (.A(net19),
    .X(data_out[7]));
 sky130_fd_sc_hd__clkbuf_4 output20 (.A(net20),
    .X(empty));
 sky130_fd_sc_hd__clkbuf_4 output21 (.A(net21),
    .X(error));
 sky130_fd_sc_hd__clkbuf_4 output22 (.A(net22),
    .X(full));
 sky130_fd_sc_hd__buf_2 max_cap23 (.A(_0217_),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_2 wire24 (.A(_0203_),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_2 wire25 (.A(_0202_),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_2 wire26 (.A(net165),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_2 wire27 (.A(net166),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\fifo[0][0] ),
    .X(net28));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\fifo[0][6] ),
    .X(net29));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\fifo[0][4] ),
    .X(net30));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\fifo[0][1] ),
    .X(net31));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\fifo[0][7] ),
    .X(net32));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\fifo[0][5] ),
    .X(net33));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\fifo[3][4] ),
    .X(net34));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\fifo[3][0] ),
    .X(net35));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\fifo[4][5] ),
    .X(net36));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\fifo[14][4] ),
    .X(net37));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\fifo[8][4] ),
    .X(net38));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\fifo[9][4] ),
    .X(net39));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\fifo[9][7] ),
    .X(net40));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\fifo[13][4] ),
    .X(net41));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\fifo[0][2] ),
    .X(net42));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\fifo[6][7] ),
    .X(net43));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\fifo[15][0] ),
    .X(net44));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\fifo[9][0] ),
    .X(net45));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\fifo[0][3] ),
    .X(net46));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\fifo[8][7] ),
    .X(net47));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\fifo[4][4] ),
    .X(net48));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\fifo[12][5] ),
    .X(net49));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\fifo[7][0] ),
    .X(net50));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\fifo[9][5] ),
    .X(net51));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\fifo[15][4] ),
    .X(net52));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\fifo[10][4] ),
    .X(net53));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\fifo[1][7] ),
    .X(net54));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\fifo[1][5] ),
    .X(net55));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\fifo[8][0] ),
    .X(net56));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\fifo[8][2] ),
    .X(net57));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\fifo[12][1] ),
    .X(net58));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\fifo[4][0] ),
    .X(net59));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\fifo[2][0] ),
    .X(net60));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\fifo[9][6] ),
    .X(net61));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\fifo[12][7] ),
    .X(net62));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(\fifo[15][5] ),
    .X(net63));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\fifo[4][6] ),
    .X(net64));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\fifo[14][0] ),
    .X(net65));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\fifo[2][7] ),
    .X(net66));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(\fifo[2][3] ),
    .X(net67));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\fifo[6][5] ),
    .X(net68));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\fifo[2][5] ),
    .X(net69));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\fifo[7][7] ),
    .X(net70));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(\fifo[3][6] ),
    .X(net71));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\fifo[11][5] ),
    .X(net72));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\fifo[8][5] ),
    .X(net73));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\fifo[6][3] ),
    .X(net74));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\fifo[6][0] ),
    .X(net75));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\fifo[10][1] ),
    .X(net76));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(\fifo[9][3] ),
    .X(net77));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\fifo[2][6] ),
    .X(net78));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(\fifo[8][1] ),
    .X(net79));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\fifo[6][4] ),
    .X(net80));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(\fifo[5][2] ),
    .X(net81));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\fifo[5][1] ),
    .X(net82));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(\fifo[12][2] ),
    .X(net83));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\fifo[6][2] ),
    .X(net84));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(\fifo[5][7] ),
    .X(net85));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(\fifo[15][1] ),
    .X(net86));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(\fifo[5][0] ),
    .X(net87));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\fifo[4][1] ),
    .X(net88));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(\fifo[1][2] ),
    .X(net89));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(\fifo[9][2] ),
    .X(net90));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(\fifo[14][1] ),
    .X(net91));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(\fifo[13][7] ),
    .X(net92));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(\fifo[13][5] ),
    .X(net93));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(\fifo[6][1] ),
    .X(net94));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(\fifo[8][3] ),
    .X(net95));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(\fifo[12][4] ),
    .X(net96));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(\fifo[1][1] ),
    .X(net97));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(\fifo[3][5] ),
    .X(net98));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(\fifo[7][5] ),
    .X(net99));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(\fifo[7][4] ),
    .X(net100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(\fifo[14][2] ),
    .X(net101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(\fifo[7][6] ),
    .X(net102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(\fifo[2][1] ),
    .X(net103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(\fifo[10][0] ),
    .X(net104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(\fifo[4][7] ),
    .X(net105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(\fifo[13][0] ),
    .X(net106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(\fifo[2][4] ),
    .X(net107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\fifo[14][5] ),
    .X(net108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(\fifo[11][0] ),
    .X(net109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(\fifo[9][1] ),
    .X(net110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(\fifo[5][4] ),
    .X(net111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\fifo[14][7] ),
    .X(net112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(\fifo[12][3] ),
    .X(net113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(\fifo[10][7] ),
    .X(net114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(\fifo[4][2] ),
    .X(net115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(\fifo[14][3] ),
    .X(net116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(\fifo[1][6] ),
    .X(net117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(\fifo[14][6] ),
    .X(net118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(\fifo[3][7] ),
    .X(net119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(\fifo[3][2] ),
    .X(net120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(\fifo[11][1] ),
    .X(net121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(\fifo[1][3] ),
    .X(net122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(\fifo[5][5] ),
    .X(net123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(\fifo[13][3] ),
    .X(net124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(\fifo[1][4] ),
    .X(net125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(\fifo[13][2] ),
    .X(net126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(\fifo[11][6] ),
    .X(net127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(\fifo[11][3] ),
    .X(net128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(\fifo[12][6] ),
    .X(net129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(\fifo[8][6] ),
    .X(net130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(\fifo[7][3] ),
    .X(net131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(\fifo[5][3] ),
    .X(net132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(\fifo[10][6] ),
    .X(net133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(\fifo[3][3] ),
    .X(net134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(\fifo[2][2] ),
    .X(net135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(\fifo[11][7] ),
    .X(net136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(\fifo[10][5] ),
    .X(net137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(\fifo[11][4] ),
    .X(net138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(\fifo[5][6] ),
    .X(net139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(\fifo[4][3] ),
    .X(net140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(\fifo[7][1] ),
    .X(net141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(\fifo[1][0] ),
    .X(net142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(\fifo[6][6] ),
    .X(net143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(\fifo[13][1] ),
    .X(net144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(\fifo[15][2] ),
    .X(net145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(\fifo[10][3] ),
    .X(net146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(\fifo[11][2] ),
    .X(net147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(\fifo[15][6] ),
    .X(net148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(\fifo[13][6] ),
    .X(net149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(\fifo[15][7] ),
    .X(net150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(\fifo[12][0] ),
    .X(net151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(\fifo[3][1] ),
    .X(net152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(\fifo[7][2] ),
    .X(net153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(\tail[4] ),
    .X(net154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(\fifo[10][2] ),
    .X(net155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(\head[4] ),
    .X(net156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(\fifo[15][3] ),
    .X(net157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(\head[3] ),
    .X(net158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(net17),
    .X(net159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(\head[1] ),
    .X(net160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(\head[2] ),
    .X(net161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(net14),
    .X(net162));
 sky130_fd_sc_hd__dlymetal6s2s_1 max_cap1 (.A(_0203_),
    .X(net163));
 sky130_fd_sc_hd__dlymetal6s2s_1 max_cap2 (.A(_0202_),
    .X(net164));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire3 (.A(_0200_),
    .X(net165));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire4 (.A(_0198_),
    .X(net166));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_31 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_107 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_59 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_330 ();
endmodule
